magic
tech scmos
timestamp 1732873084
<< nwell >>
rect 87 183 147 214
rect 93 116 153 147
rect 193 106 253 210
rect 388 204 448 235
rect 394 137 454 168
rect 494 127 554 231
rect 785 221 891 223
rect 915 221 985 223
rect 785 163 985 221
rect 1046 163 1076 223
rect 889 161 920 163
rect 191 104 253 106
rect 492 125 554 127
rect 191 80 251 104
rect 492 101 552 125
rect 492 96 554 101
rect -214 77 -108 79
rect -84 77 -14 79
rect -214 19 -14 77
rect 191 75 253 80
rect -110 17 -79 19
rect 193 10 253 75
rect 494 31 554 96
rect 781 57 812 117
rect 848 63 879 123
rect -218 -87 -187 -27
rect -151 -81 -120 -21
rect 177 -27 243 -6
rect 134 -111 159 -59
rect 176 -77 243 -27
rect 572 -32 585 -31
rect 492 -100 614 -32
rect 775 -75 881 -73
rect 905 -75 975 -73
rect 134 -112 152 -111
rect 492 -126 573 -100
rect 775 -133 975 -75
rect 1057 -133 1087 -73
rect 879 -135 910 -133
rect -111 -233 -51 -202
rect -105 -300 -45 -269
rect -5 -310 55 -206
rect 140 -243 219 -185
rect 771 -239 802 -179
rect 838 -233 869 -173
rect -7 -312 55 -310
rect -7 -336 53 -312
rect -7 -341 55 -336
rect -5 -406 55 -341
rect 154 -425 181 -373
rect 196 -392 266 -332
rect 504 -364 653 -363
rect 504 -435 688 -364
rect 849 -408 955 -406
rect 979 -408 1049 -406
rect -132 -446 -26 -444
rect -2 -446 68 -444
rect -132 -504 68 -446
rect 504 -499 599 -435
rect 849 -466 1049 -408
rect 1124 -466 1154 -406
rect 953 -468 984 -466
rect -28 -506 3 -504
rect -136 -610 -105 -550
rect -69 -604 -38 -544
rect 162 -557 241 -499
rect 845 -572 876 -512
rect 912 -566 943 -506
rect -112 -725 -6 -723
rect 18 -725 88 -723
rect -112 -783 88 -725
rect 221 -765 254 -764
rect -8 -785 23 -783
rect -116 -889 -85 -829
rect -49 -883 -18 -823
rect 155 -858 182 -802
rect 198 -820 254 -765
rect 198 -821 225 -820
rect 500 -844 696 -669
rect 842 -836 948 -834
rect 972 -836 1042 -834
rect 842 -894 1042 -836
rect 1124 -894 1154 -834
rect 946 -896 977 -894
rect 162 -986 241 -928
rect 838 -1000 869 -940
rect 905 -994 936 -934
rect -105 -1124 -45 -1059
rect -105 -1129 -43 -1124
rect -103 -1153 -43 -1129
rect -105 -1155 -43 -1153
rect -105 -1259 -45 -1155
rect 493 -1159 701 -1144
rect -5 -1196 55 -1165
rect 1 -1263 61 -1232
rect 224 -1294 257 -1293
rect -114 -1335 -8 -1333
rect 16 -1335 86 -1333
rect -114 -1393 86 -1335
rect 158 -1387 185 -1331
rect 201 -1349 257 -1294
rect 201 -1350 228 -1349
rect 493 -1362 700 -1159
rect 735 -1268 841 -1266
rect 865 -1268 935 -1266
rect 735 -1326 935 -1268
rect 1017 -1326 1047 -1266
rect 839 -1328 870 -1326
rect -10 -1395 21 -1393
rect 731 -1432 762 -1372
rect 798 -1426 829 -1366
rect -118 -1499 -87 -1439
rect -51 -1493 -20 -1433
rect 165 -1515 244 -1457
rect 63 -1664 123 -1599
rect 63 -1669 125 -1664
rect 65 -1693 125 -1669
rect 63 -1695 125 -1693
rect 63 -1799 123 -1695
rect 163 -1736 223 -1705
rect 169 -1803 229 -1772
<< ntransistor >>
rect 329 220 349 222
rect 28 199 48 201
rect 329 160 349 162
rect 28 139 48 141
rect 330 115 350 117
rect 396 109 416 111
rect 29 94 49 96
rect 95 88 115 90
rect 330 86 350 88
rect 397 86 417 88
rect 29 65 49 67
rect 397 69 417 71
rect 96 65 116 67
rect 96 48 116 50
rect 397 47 417 49
rect -94 -79 -92 -59
rect 96 26 116 28
rect -71 -78 -69 -58
rect -54 -78 -52 -58
rect -32 -78 -30 -58
rect 905 65 907 85
rect 928 66 930 86
rect 945 66 947 86
rect 967 66 969 86
rect 1058 66 1060 86
rect 794 -2 796 18
rect 854 -2 856 18
rect 899 -1 901 19
rect 928 -1 930 19
rect -205 -146 -203 -126
rect -145 -146 -143 -126
rect -100 -145 -98 -125
rect -71 -145 -69 -125
rect 189 -113 191 -94
rect 219 -113 221 -94
rect 715 -43 717 -24
rect 745 -43 747 -24
rect 671 -77 673 -58
rect 145 -147 147 -128
rect -170 -217 -150 -215
rect 510 -251 512 -211
rect 527 -251 529 -211
rect 558 -250 560 -230
rect 600 -247 602 -227
rect -170 -277 -150 -275
rect 151 -309 153 -269
rect 170 -309 172 -269
rect 205 -282 207 -262
rect 700 -255 702 -236
rect 730 -255 732 -236
rect 895 -231 897 -211
rect 656 -289 658 -270
rect 918 -230 920 -210
rect 935 -230 937 -210
rect 957 -230 959 -210
rect 1069 -230 1071 -210
rect 784 -298 786 -278
rect 844 -298 846 -278
rect 889 -297 891 -277
rect 918 -297 920 -277
rect -169 -322 -149 -320
rect -103 -328 -83 -326
rect -169 -351 -149 -349
rect -102 -351 -82 -349
rect -102 -368 -82 -366
rect -102 -390 -82 -388
rect 211 -427 213 -408
rect 241 -427 243 -408
rect 167 -461 169 -442
rect -12 -602 -10 -582
rect 11 -601 13 -581
rect 28 -601 30 -581
rect 50 -601 52 -581
rect 668 -479 670 -459
rect 776 -511 778 -492
rect 806 -511 808 -492
rect 732 -545 734 -526
rect 173 -623 175 -583
rect 192 -623 194 -583
rect 227 -596 229 -576
rect 515 -630 517 -570
rect 527 -630 529 -570
rect 546 -600 548 -570
rect 564 -630 566 -570
rect 583 -590 585 -570
rect 969 -564 971 -544
rect 992 -563 994 -543
rect 1009 -563 1011 -543
rect 1031 -563 1033 -543
rect 1136 -563 1138 -543
rect 858 -631 860 -611
rect 918 -631 920 -611
rect 963 -630 965 -610
rect 992 -630 994 -610
rect -123 -669 -121 -649
rect -63 -669 -61 -649
rect -18 -668 -16 -648
rect 11 -668 13 -648
rect 8 -881 10 -861
rect 31 -880 33 -860
rect 48 -880 50 -860
rect 70 -880 72 -860
rect 211 -856 213 -837
rect 241 -856 243 -837
rect 167 -890 169 -871
rect -103 -948 -101 -928
rect -43 -948 -41 -928
rect 2 -947 4 -927
rect 31 -947 33 -927
rect 173 -1052 175 -1012
rect 192 -1052 194 -1012
rect 227 -1025 229 -1005
rect 32 -1077 52 -1075
rect 514 -1088 516 -1008
rect 532 -1089 534 -1009
rect 550 -1088 552 -1048
rect 568 -1089 570 -1009
rect 587 -1088 589 -1062
rect 606 -1088 608 -1008
rect 767 -1028 769 -1009
rect 797 -1028 799 -1009
rect 962 -992 964 -972
rect 985 -991 987 -971
rect 1002 -991 1004 -971
rect 1024 -991 1026 -971
rect 1136 -991 1138 -971
rect 723 -1062 725 -1043
rect 851 -1059 853 -1039
rect 911 -1059 913 -1039
rect 956 -1058 958 -1038
rect 985 -1058 987 -1038
rect 624 -1088 626 -1068
rect 657 -1088 659 -1068
rect 32 -1099 52 -1097
rect 32 -1116 52 -1114
rect 99 -1116 119 -1114
rect 33 -1139 53 -1137
rect 99 -1145 119 -1143
rect 100 -1190 120 -1188
rect 100 -1250 120 -1248
rect 6 -1491 8 -1471
rect 214 -1385 216 -1366
rect 244 -1385 246 -1366
rect 170 -1419 172 -1400
rect 29 -1490 31 -1470
rect 46 -1490 48 -1470
rect 68 -1490 70 -1470
rect -105 -1558 -103 -1538
rect -45 -1558 -43 -1538
rect 0 -1557 2 -1537
rect 29 -1557 31 -1537
rect 176 -1581 178 -1541
rect 195 -1581 197 -1541
rect 230 -1554 232 -1534
rect 200 -1617 220 -1615
rect 504 -1632 506 -1532
rect 523 -1632 525 -1532
rect 541 -1632 543 -1582
rect 559 -1632 561 -1532
rect 576 -1632 578 -1599
rect 594 -1632 596 -1532
rect 612 -1632 614 -1607
rect 631 -1632 633 -1532
rect 855 -1424 857 -1404
rect 878 -1423 880 -1403
rect 895 -1423 897 -1403
rect 917 -1423 919 -1403
rect 1029 -1423 1031 -1403
rect 744 -1491 746 -1471
rect 804 -1491 806 -1471
rect 849 -1490 851 -1470
rect 878 -1490 880 -1470
rect 650 -1632 652 -1612
rect 686 -1632 688 -1612
rect 200 -1639 220 -1637
rect 200 -1656 220 -1654
rect 267 -1656 287 -1654
rect 201 -1679 221 -1677
rect 267 -1685 287 -1683
rect 268 -1730 288 -1728
rect 268 -1790 288 -1788
<< ptransistor >>
rect 400 220 439 222
rect 505 216 545 218
rect 99 199 138 201
rect 204 195 244 197
rect 798 174 800 214
rect 850 174 852 214
rect 505 164 545 166
rect 406 153 445 155
rect 204 143 244 145
rect 105 132 144 134
rect 902 172 904 212
rect 928 173 930 214
rect 945 174 947 214
rect 967 174 969 214
rect 1058 174 1060 214
rect 503 112 543 114
rect 202 91 242 93
rect 504 86 545 88
rect -201 30 -199 70
rect -149 30 -147 70
rect -97 28 -95 68
rect -71 29 -69 70
rect -54 30 -52 70
rect -32 30 -30 70
rect 505 69 545 71
rect 794 69 796 108
rect 203 65 244 67
rect 204 48 244 50
rect 505 47 545 49
rect -205 -75 -203 -36
rect -138 -69 -136 -30
rect 204 26 244 28
rect 145 -105 147 -65
rect 189 -71 191 -31
rect 219 -71 221 -31
rect 671 -35 673 5
rect 715 -1 717 39
rect 745 -1 747 39
rect 861 75 863 114
rect 510 -120 512 -40
rect 527 -120 529 -40
rect 558 -120 560 -40
rect 600 -82 602 -42
rect -99 -217 -60 -215
rect 6 -221 46 -219
rect 151 -237 153 -197
rect 170 -237 172 -197
rect 205 -237 207 -197
rect 788 -122 790 -82
rect 840 -122 842 -82
rect 892 -124 894 -84
rect 918 -123 920 -82
rect 935 -122 937 -82
rect 957 -122 959 -82
rect 1069 -122 1071 -82
rect 656 -247 658 -207
rect 700 -213 702 -173
rect 730 -213 732 -173
rect 784 -227 786 -188
rect 6 -273 46 -271
rect -93 -284 -54 -282
rect 851 -221 853 -182
rect 4 -325 44 -323
rect 5 -351 46 -349
rect 6 -368 46 -366
rect 6 -390 46 -388
rect 167 -419 169 -379
rect 211 -385 213 -345
rect 241 -385 243 -345
rect -119 -493 -117 -453
rect -67 -493 -65 -453
rect -15 -495 -13 -455
rect 11 -494 13 -453
rect 28 -493 30 -453
rect 50 -493 52 -453
rect 515 -491 517 -371
rect 527 -491 529 -371
rect -123 -598 -121 -559
rect -56 -592 -54 -553
rect 173 -551 175 -511
rect 192 -551 194 -511
rect 227 -551 229 -511
rect 546 -492 548 -372
rect 564 -432 566 -372
rect 583 -492 585 -372
rect 668 -423 670 -383
rect 732 -503 734 -463
rect 776 -469 778 -429
rect 806 -469 808 -429
rect 862 -455 864 -415
rect 914 -455 916 -415
rect 966 -457 968 -417
rect 992 -456 994 -415
rect 1009 -455 1011 -415
rect 1031 -455 1033 -415
rect 1136 -455 1138 -415
rect 858 -560 860 -521
rect 925 -554 927 -515
rect -99 -772 -97 -732
rect -47 -772 -45 -732
rect 5 -774 7 -734
rect 31 -773 33 -732
rect 48 -772 50 -732
rect 70 -772 72 -732
rect -103 -877 -101 -838
rect -36 -871 -34 -832
rect 167 -848 169 -808
rect 211 -814 213 -774
rect 241 -814 243 -774
rect 514 -838 516 -678
rect 532 -838 534 -678
rect 550 -838 552 -678
rect 568 -758 570 -678
rect 173 -980 175 -940
rect 192 -980 194 -940
rect 227 -980 229 -940
rect -96 -1077 -56 -1075
rect 587 -837 589 -677
rect 606 -731 608 -677
rect 624 -836 626 -676
rect 657 -717 659 -677
rect 855 -883 857 -843
rect 907 -883 909 -843
rect 959 -885 961 -845
rect 985 -884 987 -843
rect 1002 -883 1004 -843
rect 1024 -883 1026 -843
rect 1136 -883 1138 -843
rect 723 -1020 725 -980
rect 767 -986 769 -946
rect 797 -986 799 -946
rect 851 -988 853 -949
rect 918 -982 920 -943
rect -96 -1099 -56 -1097
rect -96 -1116 -55 -1114
rect -94 -1142 -54 -1140
rect 4 -1183 43 -1181
rect -96 -1194 -56 -1192
rect -96 -1246 -56 -1244
rect 10 -1250 49 -1248
rect -101 -1382 -99 -1342
rect -49 -1382 -47 -1342
rect 3 -1384 5 -1344
rect 29 -1383 31 -1342
rect 46 -1382 48 -1342
rect 68 -1382 70 -1342
rect 170 -1377 172 -1337
rect 214 -1343 216 -1303
rect 244 -1343 246 -1303
rect 504 -1355 506 -1155
rect 523 -1355 525 -1155
rect 541 -1355 543 -1155
rect 559 -1255 561 -1155
rect -105 -1487 -103 -1448
rect -38 -1481 -36 -1442
rect 176 -1509 178 -1469
rect 195 -1509 197 -1469
rect 230 -1509 232 -1469
rect 72 -1617 112 -1615
rect 576 -1355 578 -1155
rect 594 -1221 596 -1155
rect 612 -1355 614 -1155
rect 631 -1205 633 -1155
rect 650 -1355 652 -1155
rect 686 -1209 688 -1169
rect 748 -1315 750 -1275
rect 800 -1315 802 -1275
rect 852 -1317 854 -1277
rect 878 -1316 880 -1275
rect 895 -1315 897 -1275
rect 917 -1315 919 -1275
rect 1029 -1315 1031 -1275
rect 744 -1420 746 -1381
rect 811 -1414 813 -1375
rect 72 -1639 112 -1637
rect 72 -1656 113 -1654
rect 74 -1682 114 -1680
rect 172 -1723 211 -1721
rect 72 -1734 112 -1732
rect 72 -1786 112 -1784
rect 178 -1790 217 -1788
<< ndiffusion >>
rect 329 222 349 223
rect 329 219 349 220
rect 28 201 48 202
rect 28 198 48 199
rect 329 162 349 163
rect 329 159 349 160
rect 28 141 48 142
rect 28 138 48 139
rect 330 117 350 118
rect 330 114 350 115
rect 396 111 416 112
rect 396 108 416 109
rect 29 96 49 97
rect 29 93 49 94
rect 95 90 115 91
rect 95 87 115 88
rect 330 88 350 89
rect 397 88 417 89
rect 330 85 350 86
rect 397 85 417 86
rect 29 67 49 68
rect 96 67 116 68
rect 397 71 417 72
rect 397 68 417 69
rect 29 64 49 65
rect 96 64 116 65
rect 96 50 116 51
rect 397 49 417 50
rect 96 47 116 48
rect 397 46 417 47
rect -95 -79 -94 -59
rect -92 -79 -91 -59
rect 96 28 116 29
rect 96 25 116 26
rect -72 -78 -71 -58
rect -69 -78 -68 -58
rect -55 -78 -54 -58
rect -52 -78 -51 -58
rect -33 -78 -32 -58
rect -30 -78 -29 -58
rect 904 65 905 85
rect 907 65 908 85
rect 927 66 928 86
rect 930 66 931 86
rect 944 66 945 86
rect 947 66 948 86
rect 966 66 967 86
rect 969 66 970 86
rect 1057 66 1058 86
rect 1060 66 1061 86
rect 793 -2 794 18
rect 796 -2 797 18
rect 853 -2 854 18
rect 856 -2 857 18
rect 898 -1 899 19
rect 901 -1 902 19
rect 927 -1 928 19
rect 930 -1 931 19
rect -206 -146 -205 -126
rect -203 -146 -202 -126
rect -146 -146 -145 -126
rect -143 -146 -142 -126
rect -101 -145 -100 -125
rect -98 -145 -97 -125
rect -72 -145 -71 -125
rect -69 -145 -68 -125
rect 188 -113 189 -94
rect 191 -113 192 -94
rect 218 -113 219 -94
rect 221 -113 222 -94
rect 714 -43 715 -24
rect 717 -43 718 -24
rect 744 -43 745 -24
rect 747 -43 748 -24
rect 670 -77 671 -58
rect 673 -77 674 -58
rect 144 -147 145 -128
rect 147 -147 148 -128
rect -170 -215 -150 -214
rect -170 -218 -150 -217
rect -170 -275 -150 -274
rect 509 -251 510 -211
rect 512 -251 513 -211
rect 526 -251 527 -211
rect 529 -251 530 -211
rect 557 -250 558 -230
rect 560 -250 561 -230
rect 599 -247 600 -227
rect 602 -247 603 -227
rect -170 -278 -150 -277
rect 150 -309 151 -269
rect 153 -309 154 -269
rect 169 -309 170 -269
rect 172 -309 173 -269
rect 204 -282 205 -262
rect 207 -282 208 -262
rect 699 -255 700 -236
rect 702 -255 703 -236
rect 729 -255 730 -236
rect 732 -255 733 -236
rect 894 -231 895 -211
rect 897 -231 898 -211
rect 655 -289 656 -270
rect 658 -289 659 -270
rect 917 -230 918 -210
rect 920 -230 921 -210
rect 934 -230 935 -210
rect 937 -230 938 -210
rect 956 -230 957 -210
rect 959 -230 960 -210
rect 1068 -230 1069 -210
rect 1071 -230 1072 -210
rect 783 -298 784 -278
rect 786 -298 787 -278
rect 843 -298 844 -278
rect 846 -298 847 -278
rect 888 -297 889 -277
rect 891 -297 892 -277
rect 917 -297 918 -277
rect 920 -297 921 -277
rect -169 -320 -149 -319
rect -169 -323 -149 -322
rect -103 -326 -83 -325
rect -103 -329 -83 -328
rect -169 -349 -149 -348
rect -102 -349 -82 -348
rect -169 -352 -149 -351
rect -102 -352 -82 -351
rect -102 -366 -82 -365
rect -102 -369 -82 -368
rect -102 -388 -82 -387
rect -102 -391 -82 -390
rect 210 -427 211 -408
rect 213 -427 214 -408
rect 240 -427 241 -408
rect 243 -427 244 -408
rect 166 -461 167 -442
rect 169 -461 170 -442
rect -13 -602 -12 -582
rect -10 -602 -9 -582
rect 10 -601 11 -581
rect 13 -601 14 -581
rect 27 -601 28 -581
rect 30 -601 31 -581
rect 49 -601 50 -581
rect 52 -601 53 -581
rect 667 -479 668 -459
rect 670 -479 671 -459
rect 775 -511 776 -492
rect 778 -511 779 -492
rect 805 -511 806 -492
rect 808 -511 809 -492
rect 731 -545 732 -526
rect 734 -545 735 -526
rect 172 -623 173 -583
rect 175 -623 176 -583
rect 191 -623 192 -583
rect 194 -623 195 -583
rect 226 -596 227 -576
rect 229 -596 230 -576
rect 514 -630 515 -570
rect 517 -630 527 -570
rect 529 -630 530 -570
rect 545 -600 546 -570
rect 548 -600 549 -570
rect 563 -630 564 -570
rect 566 -630 567 -570
rect 582 -590 583 -570
rect 585 -590 586 -570
rect 968 -564 969 -544
rect 971 -564 972 -544
rect 991 -563 992 -543
rect 994 -563 995 -543
rect 1008 -563 1009 -543
rect 1011 -563 1012 -543
rect 1030 -563 1031 -543
rect 1033 -563 1034 -543
rect 1135 -563 1136 -543
rect 1138 -563 1139 -543
rect 857 -631 858 -611
rect 860 -631 861 -611
rect 917 -631 918 -611
rect 920 -631 921 -611
rect 962 -630 963 -610
rect 965 -630 966 -610
rect 991 -630 992 -610
rect 994 -630 995 -610
rect -124 -669 -123 -649
rect -121 -669 -120 -649
rect -64 -669 -63 -649
rect -61 -669 -60 -649
rect -19 -668 -18 -648
rect -16 -668 -15 -648
rect 10 -668 11 -648
rect 13 -668 14 -648
rect 7 -881 8 -861
rect 10 -881 11 -861
rect 30 -880 31 -860
rect 33 -880 34 -860
rect 47 -880 48 -860
rect 50 -880 51 -860
rect 69 -880 70 -860
rect 72 -880 73 -860
rect 210 -856 211 -837
rect 213 -856 214 -837
rect 240 -856 241 -837
rect 243 -856 244 -837
rect 166 -890 167 -871
rect 169 -890 170 -871
rect -104 -948 -103 -928
rect -101 -948 -100 -928
rect -44 -948 -43 -928
rect -41 -948 -40 -928
rect 1 -947 2 -927
rect 4 -947 5 -927
rect 30 -947 31 -927
rect 33 -947 34 -927
rect 172 -1052 173 -1012
rect 175 -1052 176 -1012
rect 191 -1052 192 -1012
rect 194 -1052 195 -1012
rect 226 -1025 227 -1005
rect 229 -1025 230 -1005
rect 32 -1075 52 -1074
rect 32 -1078 52 -1077
rect 513 -1088 514 -1008
rect 516 -1088 517 -1008
rect 531 -1089 532 -1009
rect 534 -1089 535 -1009
rect 549 -1088 550 -1048
rect 552 -1088 553 -1048
rect 567 -1089 568 -1009
rect 570 -1089 571 -1009
rect 586 -1088 587 -1062
rect 589 -1088 590 -1062
rect 605 -1088 606 -1008
rect 608 -1088 609 -1008
rect 766 -1028 767 -1009
rect 769 -1028 770 -1009
rect 796 -1028 797 -1009
rect 799 -1028 800 -1009
rect 961 -992 962 -972
rect 964 -992 965 -972
rect 984 -991 985 -971
rect 987 -991 988 -971
rect 1001 -991 1002 -971
rect 1004 -991 1005 -971
rect 1023 -991 1024 -971
rect 1026 -991 1027 -971
rect 1135 -991 1136 -971
rect 1138 -991 1139 -971
rect 722 -1062 723 -1043
rect 725 -1062 726 -1043
rect 850 -1059 851 -1039
rect 853 -1059 854 -1039
rect 910 -1059 911 -1039
rect 913 -1059 914 -1039
rect 955 -1058 956 -1038
rect 958 -1058 959 -1038
rect 984 -1058 985 -1038
rect 987 -1058 988 -1038
rect 623 -1088 624 -1068
rect 626 -1088 627 -1068
rect 656 -1088 657 -1068
rect 659 -1088 660 -1068
rect 32 -1097 52 -1096
rect 32 -1100 52 -1099
rect 32 -1114 52 -1113
rect 99 -1114 119 -1113
rect 32 -1117 52 -1116
rect 99 -1117 119 -1116
rect 33 -1137 53 -1136
rect 33 -1140 53 -1139
rect 99 -1143 119 -1142
rect 99 -1146 119 -1145
rect 100 -1188 120 -1187
rect 100 -1191 120 -1190
rect 100 -1248 120 -1247
rect 100 -1251 120 -1250
rect 5 -1491 6 -1471
rect 8 -1491 9 -1471
rect 213 -1385 214 -1366
rect 216 -1385 217 -1366
rect 243 -1385 244 -1366
rect 246 -1385 247 -1366
rect 169 -1419 170 -1400
rect 172 -1419 173 -1400
rect 28 -1490 29 -1470
rect 31 -1490 32 -1470
rect 45 -1490 46 -1470
rect 48 -1490 49 -1470
rect 67 -1490 68 -1470
rect 70 -1490 71 -1470
rect -106 -1558 -105 -1538
rect -103 -1558 -102 -1538
rect -46 -1558 -45 -1538
rect -43 -1558 -42 -1538
rect -1 -1557 0 -1537
rect 2 -1557 3 -1537
rect 28 -1557 29 -1537
rect 31 -1557 32 -1537
rect 175 -1581 176 -1541
rect 178 -1581 179 -1541
rect 194 -1581 195 -1541
rect 197 -1581 198 -1541
rect 229 -1554 230 -1534
rect 232 -1554 233 -1534
rect 200 -1615 220 -1614
rect 200 -1618 220 -1617
rect 503 -1632 504 -1532
rect 506 -1632 507 -1532
rect 522 -1632 523 -1532
rect 525 -1632 526 -1532
rect 540 -1632 541 -1582
rect 543 -1632 544 -1582
rect 558 -1632 559 -1532
rect 561 -1632 562 -1532
rect 575 -1632 576 -1599
rect 578 -1632 579 -1599
rect 593 -1632 594 -1532
rect 596 -1632 597 -1532
rect 611 -1632 612 -1607
rect 614 -1632 615 -1607
rect 630 -1632 631 -1532
rect 633 -1632 634 -1532
rect 854 -1424 855 -1404
rect 857 -1424 858 -1404
rect 877 -1423 878 -1403
rect 880 -1423 881 -1403
rect 894 -1423 895 -1403
rect 897 -1423 898 -1403
rect 916 -1423 917 -1403
rect 919 -1423 920 -1403
rect 1028 -1423 1029 -1403
rect 1031 -1423 1032 -1403
rect 743 -1491 744 -1471
rect 746 -1491 747 -1471
rect 803 -1491 804 -1471
rect 806 -1491 807 -1471
rect 848 -1490 849 -1470
rect 851 -1490 852 -1470
rect 877 -1490 878 -1470
rect 880 -1490 881 -1470
rect 649 -1632 650 -1612
rect 652 -1632 653 -1612
rect 685 -1632 686 -1612
rect 688 -1632 689 -1612
rect 200 -1637 220 -1636
rect 200 -1640 220 -1639
rect 200 -1654 220 -1653
rect 267 -1654 287 -1653
rect 200 -1657 220 -1656
rect 267 -1657 287 -1656
rect 201 -1677 221 -1676
rect 201 -1680 221 -1679
rect 267 -1683 287 -1682
rect 267 -1686 287 -1685
rect 268 -1728 288 -1727
rect 268 -1731 288 -1730
rect 268 -1788 288 -1787
rect 268 -1791 288 -1790
<< pdiffusion >>
rect 400 222 439 223
rect 400 219 439 220
rect 505 218 545 219
rect 505 215 545 216
rect 99 201 138 202
rect 99 198 138 199
rect 204 197 244 198
rect 204 194 244 195
rect 797 174 798 214
rect 800 174 801 214
rect 849 174 850 214
rect 852 174 853 214
rect 505 166 545 167
rect 505 163 545 164
rect 406 155 445 156
rect 406 152 445 153
rect 204 145 244 146
rect 204 142 244 143
rect 105 134 144 135
rect 105 131 144 132
rect 901 172 902 212
rect 904 172 905 212
rect 927 173 928 214
rect 930 173 931 214
rect 944 174 945 214
rect 947 174 948 214
rect 966 174 967 214
rect 969 174 970 214
rect 1057 174 1058 214
rect 1060 174 1061 214
rect 503 114 543 115
rect 503 111 543 112
rect 202 93 242 94
rect 202 90 242 91
rect 504 88 545 89
rect 504 85 545 86
rect -202 30 -201 70
rect -199 30 -198 70
rect -150 30 -149 70
rect -147 30 -146 70
rect -98 28 -97 68
rect -95 28 -94 68
rect -72 29 -71 70
rect -69 29 -68 70
rect -55 30 -54 70
rect -52 30 -51 70
rect -33 30 -32 70
rect -30 30 -29 70
rect 505 71 545 72
rect 793 69 794 108
rect 796 69 797 108
rect 203 67 244 68
rect 203 64 244 65
rect 505 68 545 69
rect 204 50 244 51
rect 505 49 545 50
rect 204 47 244 48
rect 505 46 545 47
rect -206 -75 -205 -36
rect -203 -75 -202 -36
rect -139 -69 -138 -30
rect -136 -69 -135 -30
rect 204 28 244 29
rect 204 25 244 26
rect 144 -105 145 -65
rect 147 -105 148 -65
rect 188 -71 189 -31
rect 191 -71 192 -31
rect 218 -71 219 -31
rect 221 -71 222 -31
rect 670 -35 671 5
rect 673 -35 674 5
rect 714 -1 715 39
rect 717 -1 718 39
rect 744 -1 745 39
rect 747 -1 748 39
rect 860 75 861 114
rect 863 75 864 114
rect 509 -120 510 -40
rect 512 -120 513 -40
rect 526 -120 527 -40
rect 529 -120 530 -40
rect 557 -120 558 -40
rect 560 -120 561 -40
rect 599 -82 600 -42
rect 602 -82 603 -42
rect -99 -215 -60 -214
rect -99 -218 -60 -217
rect 6 -219 46 -218
rect 6 -222 46 -221
rect 150 -237 151 -197
rect 153 -237 154 -197
rect 169 -237 170 -197
rect 172 -237 173 -197
rect 204 -237 205 -197
rect 207 -237 208 -197
rect 787 -122 788 -82
rect 790 -122 791 -82
rect 839 -122 840 -82
rect 842 -122 843 -82
rect 891 -124 892 -84
rect 894 -124 895 -84
rect 917 -123 918 -82
rect 920 -123 921 -82
rect 934 -122 935 -82
rect 937 -122 938 -82
rect 956 -122 957 -82
rect 959 -122 960 -82
rect 1068 -122 1069 -82
rect 1071 -122 1072 -82
rect 655 -247 656 -207
rect 658 -247 659 -207
rect 699 -213 700 -173
rect 702 -213 703 -173
rect 729 -213 730 -173
rect 732 -213 733 -173
rect 783 -227 784 -188
rect 786 -227 787 -188
rect 6 -271 46 -270
rect 6 -274 46 -273
rect -93 -282 -54 -281
rect -93 -285 -54 -284
rect 850 -221 851 -182
rect 853 -221 854 -182
rect 4 -323 44 -322
rect 4 -326 44 -325
rect 5 -349 46 -348
rect 5 -352 46 -351
rect 6 -366 46 -365
rect 6 -369 46 -368
rect 6 -388 46 -387
rect 6 -391 46 -390
rect 166 -419 167 -379
rect 169 -419 170 -379
rect 210 -385 211 -345
rect 213 -385 214 -345
rect 240 -385 241 -345
rect 243 -385 244 -345
rect -120 -493 -119 -453
rect -117 -493 -116 -453
rect -68 -493 -67 -453
rect -65 -493 -64 -453
rect -16 -495 -15 -455
rect -13 -495 -12 -455
rect 10 -494 11 -453
rect 13 -494 14 -453
rect 27 -493 28 -453
rect 30 -493 31 -453
rect 49 -493 50 -453
rect 52 -493 53 -453
rect 514 -491 515 -371
rect 517 -491 520 -371
rect 524 -491 527 -371
rect 529 -491 530 -371
rect -124 -598 -123 -559
rect -121 -598 -120 -559
rect -57 -592 -56 -553
rect -54 -592 -53 -553
rect 172 -551 173 -511
rect 175 -551 176 -511
rect 191 -551 192 -511
rect 194 -551 195 -511
rect 226 -551 227 -511
rect 229 -551 230 -511
rect 545 -492 546 -372
rect 548 -492 549 -372
rect 563 -432 564 -372
rect 566 -432 567 -372
rect 582 -492 583 -372
rect 585 -492 586 -372
rect 667 -423 668 -383
rect 670 -423 671 -383
rect 731 -503 732 -463
rect 734 -503 735 -463
rect 775 -469 776 -429
rect 778 -469 779 -429
rect 805 -469 806 -429
rect 808 -469 809 -429
rect 861 -455 862 -415
rect 864 -455 865 -415
rect 913 -455 914 -415
rect 916 -455 917 -415
rect 965 -457 966 -417
rect 968 -457 969 -417
rect 991 -456 992 -415
rect 994 -456 995 -415
rect 1008 -455 1009 -415
rect 1011 -455 1012 -415
rect 1030 -455 1031 -415
rect 1033 -455 1034 -415
rect 1135 -455 1136 -415
rect 1138 -455 1139 -415
rect 857 -560 858 -521
rect 860 -560 861 -521
rect 924 -554 925 -515
rect 927 -554 928 -515
rect -100 -772 -99 -732
rect -97 -772 -96 -732
rect -48 -772 -47 -732
rect -45 -772 -44 -732
rect 4 -774 5 -734
rect 7 -774 8 -734
rect 30 -773 31 -732
rect 33 -773 34 -732
rect 47 -772 48 -732
rect 50 -772 51 -732
rect 69 -772 70 -732
rect 72 -772 73 -732
rect -104 -877 -103 -838
rect -101 -877 -100 -838
rect -37 -871 -36 -832
rect -34 -871 -33 -832
rect 166 -848 167 -808
rect 169 -848 170 -808
rect 210 -814 211 -774
rect 213 -814 214 -774
rect 240 -814 241 -774
rect 243 -814 244 -774
rect 513 -838 514 -678
rect 516 -838 517 -678
rect 531 -838 532 -678
rect 534 -838 535 -678
rect 549 -838 550 -678
rect 552 -838 553 -678
rect 567 -758 568 -678
rect 570 -758 571 -678
rect 172 -980 173 -940
rect 175 -980 176 -940
rect 191 -980 192 -940
rect 194 -980 195 -940
rect 226 -980 227 -940
rect 229 -980 230 -940
rect -96 -1075 -56 -1074
rect -96 -1078 -56 -1077
rect 586 -837 587 -677
rect 589 -837 590 -677
rect 605 -731 606 -677
rect 608 -731 609 -677
rect 623 -836 624 -676
rect 626 -836 627 -676
rect 656 -717 657 -677
rect 659 -717 660 -677
rect 854 -883 855 -843
rect 857 -883 858 -843
rect 906 -883 907 -843
rect 909 -883 910 -843
rect 958 -885 959 -845
rect 961 -885 962 -845
rect 984 -884 985 -843
rect 987 -884 988 -843
rect 1001 -883 1002 -843
rect 1004 -883 1005 -843
rect 1023 -883 1024 -843
rect 1026 -883 1027 -843
rect 1135 -883 1136 -843
rect 1138 -883 1139 -843
rect 722 -1020 723 -980
rect 725 -1020 726 -980
rect 766 -986 767 -946
rect 769 -986 770 -946
rect 796 -986 797 -946
rect 799 -986 800 -946
rect 850 -988 851 -949
rect 853 -988 854 -949
rect 917 -982 918 -943
rect 920 -982 921 -943
rect -96 -1097 -56 -1096
rect -96 -1100 -56 -1099
rect -96 -1114 -55 -1113
rect -96 -1117 -55 -1116
rect -94 -1140 -54 -1139
rect -94 -1143 -54 -1142
rect 4 -1181 43 -1180
rect 4 -1184 43 -1183
rect -96 -1192 -56 -1191
rect -96 -1195 -56 -1194
rect -96 -1244 -56 -1243
rect -96 -1247 -56 -1246
rect 10 -1248 49 -1247
rect 10 -1251 49 -1250
rect -102 -1382 -101 -1342
rect -99 -1382 -98 -1342
rect -50 -1382 -49 -1342
rect -47 -1382 -46 -1342
rect 2 -1384 3 -1344
rect 5 -1384 6 -1344
rect 28 -1383 29 -1342
rect 31 -1383 32 -1342
rect 45 -1382 46 -1342
rect 48 -1382 49 -1342
rect 67 -1382 68 -1342
rect 70 -1382 71 -1342
rect 169 -1377 170 -1337
rect 172 -1377 173 -1337
rect 213 -1343 214 -1303
rect 216 -1343 217 -1303
rect 243 -1343 244 -1303
rect 246 -1343 247 -1303
rect 503 -1355 504 -1155
rect 506 -1355 507 -1155
rect 522 -1355 523 -1155
rect 525 -1355 526 -1155
rect 540 -1355 541 -1155
rect 543 -1355 544 -1155
rect 558 -1255 559 -1155
rect 561 -1255 562 -1155
rect -106 -1487 -105 -1448
rect -103 -1487 -102 -1448
rect -39 -1481 -38 -1442
rect -36 -1481 -35 -1442
rect 175 -1509 176 -1469
rect 178 -1509 179 -1469
rect 194 -1509 195 -1469
rect 197 -1509 198 -1469
rect 229 -1509 230 -1469
rect 232 -1509 233 -1469
rect 72 -1615 112 -1614
rect 72 -1618 112 -1617
rect 575 -1355 576 -1155
rect 578 -1355 579 -1155
rect 593 -1221 594 -1155
rect 596 -1221 597 -1155
rect 611 -1355 612 -1155
rect 614 -1355 615 -1155
rect 630 -1205 631 -1155
rect 633 -1205 634 -1155
rect 649 -1355 650 -1155
rect 652 -1355 653 -1155
rect 685 -1209 686 -1169
rect 688 -1209 689 -1169
rect 747 -1315 748 -1275
rect 750 -1315 751 -1275
rect 799 -1315 800 -1275
rect 802 -1315 803 -1275
rect 851 -1317 852 -1277
rect 854 -1317 855 -1277
rect 877 -1316 878 -1275
rect 880 -1316 881 -1275
rect 894 -1315 895 -1275
rect 897 -1315 898 -1275
rect 916 -1315 917 -1275
rect 919 -1315 920 -1275
rect 1028 -1315 1029 -1275
rect 1031 -1315 1032 -1275
rect 743 -1420 744 -1381
rect 746 -1420 747 -1381
rect 810 -1414 811 -1375
rect 813 -1414 814 -1375
rect 72 -1637 112 -1636
rect 72 -1640 112 -1639
rect 72 -1654 113 -1653
rect 72 -1657 113 -1656
rect 74 -1680 114 -1679
rect 74 -1683 114 -1682
rect 172 -1721 211 -1720
rect 172 -1724 211 -1723
rect 72 -1732 112 -1731
rect 72 -1735 112 -1734
rect 72 -1784 112 -1783
rect 72 -1787 112 -1786
rect 178 -1788 217 -1787
rect 178 -1791 217 -1790
<< ndcontact >>
rect 329 223 349 227
rect 329 215 349 219
rect 28 202 48 206
rect 28 194 48 198
rect 329 163 349 167
rect 329 155 349 159
rect 28 142 48 146
rect 28 134 48 138
rect 330 118 350 122
rect 330 110 350 114
rect 396 112 416 116
rect 396 104 416 108
rect 29 97 49 101
rect 29 89 49 93
rect 95 91 115 95
rect 95 83 115 87
rect 330 89 350 93
rect 397 89 417 93
rect 330 81 350 85
rect 397 81 417 85
rect 29 68 49 72
rect 96 68 116 72
rect 397 72 417 76
rect 29 60 49 64
rect 96 60 116 64
rect 397 64 417 68
rect 96 51 116 55
rect 397 50 417 54
rect 96 43 116 47
rect 397 42 417 46
rect -99 -79 -95 -59
rect -91 -79 -87 -59
rect 96 29 116 33
rect 96 21 116 25
rect -76 -78 -72 -58
rect -68 -78 -64 -58
rect -59 -78 -55 -58
rect -51 -78 -47 -58
rect -37 -78 -33 -58
rect -29 -78 -25 -58
rect 900 65 904 85
rect 908 65 912 85
rect 923 66 927 86
rect 931 66 935 86
rect 940 66 944 86
rect 948 66 952 86
rect 962 66 966 86
rect 970 66 974 86
rect 1053 66 1057 86
rect 1061 66 1065 86
rect 789 -2 793 18
rect 797 -2 801 18
rect 849 -2 853 18
rect 857 -2 861 18
rect 894 -1 898 19
rect 902 -1 906 19
rect 923 -1 927 19
rect 931 -1 935 19
rect -210 -146 -206 -126
rect -202 -146 -198 -126
rect -150 -146 -146 -126
rect -142 -146 -138 -126
rect -105 -145 -101 -125
rect -97 -145 -93 -125
rect -76 -145 -72 -125
rect -68 -145 -64 -125
rect 184 -113 188 -94
rect 192 -113 196 -94
rect 214 -113 218 -94
rect 222 -113 226 -94
rect 710 -43 714 -24
rect 718 -43 722 -24
rect 740 -43 744 -24
rect 748 -43 752 -24
rect 666 -77 670 -58
rect 674 -77 678 -58
rect 140 -147 144 -128
rect 148 -147 152 -128
rect -170 -214 -150 -210
rect -170 -222 -150 -218
rect -170 -274 -150 -270
rect 505 -251 509 -211
rect 513 -251 517 -211
rect 522 -251 526 -211
rect 530 -251 534 -211
rect 553 -250 557 -230
rect 561 -250 565 -230
rect 595 -247 599 -227
rect 603 -247 607 -227
rect -170 -282 -150 -278
rect 146 -309 150 -269
rect 154 -309 158 -269
rect 165 -309 169 -269
rect 173 -309 177 -269
rect 200 -282 204 -262
rect 208 -282 212 -262
rect 695 -255 699 -236
rect 703 -255 707 -236
rect 725 -255 729 -236
rect 733 -255 737 -236
rect 890 -231 894 -211
rect 898 -231 902 -211
rect 651 -289 655 -270
rect 659 -289 663 -270
rect 913 -230 917 -210
rect 921 -230 925 -210
rect 930 -230 934 -210
rect 938 -230 942 -210
rect 952 -230 956 -210
rect 960 -230 964 -210
rect 1064 -230 1068 -210
rect 1072 -230 1076 -210
rect 779 -298 783 -278
rect 787 -298 791 -278
rect 839 -298 843 -278
rect 847 -298 851 -278
rect 884 -297 888 -277
rect 892 -297 896 -277
rect 913 -297 917 -277
rect 921 -297 925 -277
rect -169 -319 -149 -315
rect -169 -327 -149 -323
rect -103 -325 -83 -321
rect -103 -333 -83 -329
rect -169 -348 -149 -344
rect -102 -348 -82 -344
rect -169 -356 -149 -352
rect -102 -356 -82 -352
rect -102 -365 -82 -361
rect -102 -373 -82 -369
rect -102 -387 -82 -383
rect -102 -395 -82 -391
rect 206 -427 210 -408
rect 214 -427 218 -408
rect 236 -427 240 -408
rect 244 -427 248 -408
rect 162 -461 166 -442
rect 170 -461 174 -442
rect -17 -602 -13 -582
rect -9 -602 -5 -582
rect 6 -601 10 -581
rect 14 -601 18 -581
rect 23 -601 27 -581
rect 31 -601 35 -581
rect 45 -601 49 -581
rect 53 -601 57 -581
rect 663 -479 667 -459
rect 671 -479 675 -459
rect 771 -511 775 -492
rect 779 -511 783 -492
rect 801 -511 805 -492
rect 809 -511 813 -492
rect 727 -545 731 -526
rect 735 -545 739 -526
rect 168 -623 172 -583
rect 176 -623 180 -583
rect 187 -623 191 -583
rect 195 -623 199 -583
rect 222 -596 226 -576
rect 230 -596 234 -576
rect 510 -630 514 -570
rect 530 -630 534 -570
rect 541 -600 545 -570
rect 549 -600 553 -570
rect 559 -630 563 -570
rect 567 -630 571 -570
rect 578 -590 582 -570
rect 586 -590 590 -570
rect 964 -564 968 -544
rect 972 -564 976 -544
rect 987 -563 991 -543
rect 995 -563 999 -543
rect 1004 -563 1008 -543
rect 1012 -563 1016 -543
rect 1026 -563 1030 -543
rect 1034 -563 1038 -543
rect 1131 -563 1135 -543
rect 1139 -563 1143 -543
rect 853 -631 857 -611
rect 861 -631 865 -611
rect 913 -631 917 -611
rect 921 -631 925 -611
rect 958 -630 962 -610
rect 966 -630 970 -610
rect 987 -630 991 -610
rect 995 -630 999 -610
rect -128 -669 -124 -649
rect -120 -669 -116 -649
rect -68 -669 -64 -649
rect -60 -669 -56 -649
rect -23 -668 -19 -648
rect -15 -668 -11 -648
rect 6 -668 10 -648
rect 14 -668 18 -648
rect 3 -881 7 -861
rect 11 -881 15 -861
rect 26 -880 30 -860
rect 34 -880 38 -860
rect 43 -880 47 -860
rect 51 -880 55 -860
rect 65 -880 69 -860
rect 73 -880 77 -860
rect 206 -856 210 -837
rect 214 -856 218 -837
rect 236 -856 240 -837
rect 244 -856 248 -837
rect 162 -890 166 -871
rect 170 -890 174 -871
rect -108 -948 -104 -928
rect -100 -948 -96 -928
rect -48 -948 -44 -928
rect -40 -948 -36 -928
rect -3 -947 1 -927
rect 5 -947 9 -927
rect 26 -947 30 -927
rect 34 -947 38 -927
rect 168 -1052 172 -1012
rect 176 -1052 180 -1012
rect 187 -1052 191 -1012
rect 195 -1052 199 -1012
rect 222 -1025 226 -1005
rect 230 -1025 234 -1005
rect 32 -1074 52 -1070
rect 32 -1082 52 -1078
rect 509 -1088 513 -1008
rect 517 -1088 521 -1008
rect 527 -1089 531 -1009
rect 535 -1089 539 -1009
rect 545 -1088 549 -1048
rect 553 -1088 557 -1048
rect 563 -1089 567 -1009
rect 571 -1089 575 -1009
rect 582 -1088 586 -1062
rect 590 -1088 594 -1062
rect 601 -1088 605 -1008
rect 609 -1088 613 -1008
rect 762 -1028 766 -1009
rect 770 -1028 774 -1009
rect 792 -1028 796 -1009
rect 800 -1028 804 -1009
rect 957 -992 961 -972
rect 965 -992 969 -972
rect 980 -991 984 -971
rect 988 -991 992 -971
rect 997 -991 1001 -971
rect 1005 -991 1009 -971
rect 1019 -991 1023 -971
rect 1027 -991 1031 -971
rect 1131 -991 1135 -971
rect 1139 -991 1143 -971
rect 718 -1062 722 -1043
rect 726 -1062 730 -1043
rect 846 -1059 850 -1039
rect 854 -1059 858 -1039
rect 906 -1059 910 -1039
rect 914 -1059 918 -1039
rect 951 -1058 955 -1038
rect 959 -1058 963 -1038
rect 980 -1058 984 -1038
rect 988 -1058 992 -1038
rect 619 -1088 623 -1068
rect 627 -1088 631 -1068
rect 652 -1088 656 -1068
rect 660 -1088 664 -1068
rect 32 -1096 52 -1092
rect 32 -1104 52 -1100
rect 32 -1113 52 -1109
rect 99 -1113 119 -1109
rect 32 -1121 52 -1117
rect 99 -1121 119 -1117
rect 33 -1136 53 -1132
rect 33 -1144 53 -1140
rect 99 -1142 119 -1138
rect 99 -1150 119 -1146
rect 100 -1187 120 -1183
rect 100 -1195 120 -1191
rect 100 -1247 120 -1243
rect 100 -1255 120 -1251
rect 1 -1491 5 -1471
rect 9 -1491 13 -1471
rect 209 -1385 213 -1366
rect 217 -1385 221 -1366
rect 239 -1385 243 -1366
rect 247 -1385 251 -1366
rect 165 -1419 169 -1400
rect 173 -1419 177 -1400
rect 24 -1490 28 -1470
rect 32 -1490 36 -1470
rect 41 -1490 45 -1470
rect 49 -1490 53 -1470
rect 63 -1490 67 -1470
rect 71 -1490 75 -1470
rect -110 -1558 -106 -1538
rect -102 -1558 -98 -1538
rect -50 -1558 -46 -1538
rect -42 -1558 -38 -1538
rect -5 -1557 -1 -1537
rect 3 -1557 7 -1537
rect 24 -1557 28 -1537
rect 32 -1557 36 -1537
rect 171 -1581 175 -1541
rect 179 -1581 183 -1541
rect 190 -1581 194 -1541
rect 198 -1581 202 -1541
rect 225 -1554 229 -1534
rect 233 -1554 237 -1534
rect 200 -1614 220 -1610
rect 200 -1622 220 -1618
rect 499 -1632 503 -1532
rect 507 -1632 511 -1532
rect 518 -1632 522 -1532
rect 526 -1632 530 -1532
rect 536 -1632 540 -1582
rect 544 -1632 548 -1582
rect 554 -1632 558 -1532
rect 562 -1632 566 -1532
rect 571 -1632 575 -1599
rect 579 -1632 583 -1599
rect 589 -1632 593 -1532
rect 597 -1632 601 -1532
rect 607 -1632 611 -1607
rect 615 -1632 619 -1607
rect 626 -1632 630 -1532
rect 634 -1632 638 -1532
rect 850 -1424 854 -1404
rect 858 -1424 862 -1404
rect 873 -1423 877 -1403
rect 881 -1423 885 -1403
rect 890 -1423 894 -1403
rect 898 -1423 902 -1403
rect 912 -1423 916 -1403
rect 920 -1423 924 -1403
rect 1024 -1423 1028 -1403
rect 1032 -1423 1036 -1403
rect 739 -1491 743 -1471
rect 747 -1491 751 -1471
rect 799 -1491 803 -1471
rect 807 -1491 811 -1471
rect 844 -1490 848 -1470
rect 852 -1490 856 -1470
rect 873 -1490 877 -1470
rect 881 -1490 885 -1470
rect 645 -1632 649 -1612
rect 653 -1632 657 -1612
rect 681 -1632 685 -1612
rect 689 -1632 693 -1612
rect 200 -1636 220 -1632
rect 200 -1644 220 -1640
rect 200 -1653 220 -1649
rect 267 -1653 287 -1649
rect 200 -1661 220 -1657
rect 267 -1661 287 -1657
rect 201 -1676 221 -1672
rect 201 -1684 221 -1680
rect 267 -1682 287 -1678
rect 267 -1690 287 -1686
rect 268 -1727 288 -1723
rect 268 -1735 288 -1731
rect 268 -1787 288 -1783
rect 268 -1795 288 -1791
<< pdcontact >>
rect 400 223 439 227
rect 400 215 439 219
rect 505 219 545 223
rect 505 211 545 215
rect 99 202 138 206
rect 99 194 138 198
rect 204 198 244 202
rect 204 190 244 194
rect 793 174 797 214
rect 801 174 805 214
rect 845 174 849 214
rect 853 174 857 214
rect 505 167 545 171
rect 406 156 445 160
rect 505 159 545 163
rect 204 146 244 150
rect 406 148 445 152
rect 105 135 144 139
rect 204 138 244 142
rect 105 127 144 131
rect 897 172 901 212
rect 905 172 909 212
rect 923 173 927 214
rect 931 173 935 214
rect 940 174 944 214
rect 948 174 952 214
rect 962 174 966 214
rect 970 174 974 214
rect 1053 174 1057 214
rect 1061 174 1065 214
rect 503 115 543 119
rect 503 107 543 111
rect 202 94 242 98
rect 202 86 242 90
rect 504 89 545 93
rect 504 81 545 85
rect -206 30 -202 70
rect -198 30 -194 70
rect -154 30 -150 70
rect -146 30 -142 70
rect -102 28 -98 68
rect -94 28 -90 68
rect -76 29 -72 70
rect -68 29 -64 70
rect -59 30 -55 70
rect -51 30 -47 70
rect -37 30 -33 70
rect -29 30 -25 70
rect 203 68 244 72
rect 505 72 545 76
rect 789 69 793 108
rect 797 69 801 108
rect 505 64 545 68
rect 203 60 244 64
rect 204 51 244 55
rect 505 50 545 54
rect 204 43 244 47
rect 505 42 545 46
rect -210 -75 -206 -36
rect -202 -75 -198 -36
rect -143 -69 -139 -30
rect -135 -69 -131 -30
rect 204 29 244 33
rect 204 21 244 25
rect 140 -105 144 -65
rect 148 -105 152 -65
rect 184 -71 188 -31
rect 192 -71 196 -31
rect 214 -71 218 -31
rect 222 -71 226 -31
rect 666 -35 670 5
rect 674 -35 678 5
rect 710 -1 714 39
rect 718 -1 722 39
rect 740 -1 744 39
rect 748 -1 752 39
rect 856 75 860 114
rect 864 75 868 114
rect 505 -120 509 -40
rect 513 -120 517 -40
rect 522 -120 526 -40
rect 530 -120 534 -40
rect 553 -120 557 -40
rect 561 -120 565 -40
rect 595 -82 599 -42
rect 603 -82 607 -42
rect -99 -214 -60 -210
rect -99 -222 -60 -218
rect 6 -218 46 -214
rect 6 -226 46 -222
rect 146 -237 150 -197
rect 154 -237 158 -197
rect 165 -237 169 -197
rect 173 -237 177 -197
rect 200 -237 204 -197
rect 208 -237 212 -197
rect 6 -270 46 -266
rect 783 -122 787 -82
rect 791 -122 795 -82
rect 835 -122 839 -82
rect 843 -122 847 -82
rect 887 -124 891 -84
rect 895 -124 899 -84
rect 913 -123 917 -82
rect 921 -123 925 -82
rect 930 -122 934 -82
rect 938 -122 942 -82
rect 952 -122 956 -82
rect 960 -122 964 -82
rect 1064 -122 1068 -82
rect 1072 -122 1076 -82
rect 651 -247 655 -207
rect 659 -247 663 -207
rect 695 -213 699 -173
rect 703 -213 707 -173
rect 725 -213 729 -173
rect 733 -213 737 -173
rect 779 -227 783 -188
rect 787 -227 791 -188
rect -93 -281 -54 -277
rect 6 -278 46 -274
rect -93 -289 -54 -285
rect 846 -221 850 -182
rect 854 -221 858 -182
rect 4 -322 44 -318
rect 4 -330 44 -326
rect 5 -348 46 -344
rect 5 -356 46 -352
rect 6 -365 46 -361
rect 6 -373 46 -369
rect 6 -387 46 -383
rect 6 -395 46 -391
rect 162 -419 166 -379
rect 170 -419 174 -379
rect 206 -385 210 -345
rect 214 -385 218 -345
rect 236 -385 240 -345
rect 244 -385 248 -345
rect -124 -493 -120 -453
rect -116 -493 -112 -453
rect -72 -493 -68 -453
rect -64 -493 -60 -453
rect -20 -495 -16 -455
rect -12 -495 -8 -455
rect 6 -494 10 -453
rect 14 -494 18 -453
rect 23 -493 27 -453
rect 31 -493 35 -453
rect 45 -493 49 -453
rect 53 -493 57 -453
rect 510 -491 514 -371
rect 520 -491 524 -371
rect 530 -491 534 -371
rect -128 -598 -124 -559
rect -120 -598 -116 -559
rect -61 -592 -57 -553
rect -53 -592 -49 -553
rect 168 -551 172 -511
rect 176 -551 180 -511
rect 187 -551 191 -511
rect 195 -551 199 -511
rect 222 -551 226 -511
rect 230 -551 234 -511
rect 541 -492 545 -372
rect 549 -492 553 -372
rect 559 -432 563 -372
rect 567 -432 571 -372
rect 578 -492 582 -372
rect 586 -492 590 -372
rect 663 -423 667 -383
rect 671 -423 675 -383
rect 727 -503 731 -463
rect 735 -503 739 -463
rect 771 -469 775 -429
rect 779 -469 783 -429
rect 801 -469 805 -429
rect 809 -469 813 -429
rect 857 -455 861 -415
rect 865 -455 869 -415
rect 909 -455 913 -415
rect 917 -455 921 -415
rect 961 -457 965 -417
rect 969 -457 973 -417
rect 987 -456 991 -415
rect 995 -456 999 -415
rect 1004 -455 1008 -415
rect 1012 -455 1016 -415
rect 1026 -455 1030 -415
rect 1034 -455 1038 -415
rect 1131 -455 1135 -415
rect 1139 -455 1143 -415
rect 853 -560 857 -521
rect 861 -560 865 -521
rect 920 -554 924 -515
rect 928 -554 932 -515
rect -104 -772 -100 -732
rect -96 -772 -92 -732
rect -52 -772 -48 -732
rect -44 -772 -40 -732
rect 0 -774 4 -734
rect 8 -774 12 -734
rect 26 -773 30 -732
rect 34 -773 38 -732
rect 43 -772 47 -732
rect 51 -772 55 -732
rect 65 -772 69 -732
rect 73 -772 77 -732
rect -108 -877 -104 -838
rect -100 -877 -96 -838
rect -41 -871 -37 -832
rect -33 -871 -29 -832
rect 162 -848 166 -808
rect 170 -848 174 -808
rect 206 -814 210 -774
rect 214 -814 218 -774
rect 236 -814 240 -774
rect 244 -814 248 -774
rect 509 -838 513 -678
rect 517 -838 521 -678
rect 527 -838 531 -678
rect 535 -838 539 -678
rect 545 -838 549 -678
rect 553 -838 557 -678
rect 563 -758 567 -678
rect 571 -758 575 -678
rect 168 -980 172 -940
rect 176 -980 180 -940
rect 187 -980 191 -940
rect 195 -980 199 -940
rect 222 -980 226 -940
rect 230 -980 234 -940
rect -96 -1074 -56 -1070
rect -96 -1082 -56 -1078
rect 582 -837 586 -677
rect 590 -837 594 -677
rect 601 -731 605 -677
rect 609 -731 613 -677
rect 619 -836 623 -676
rect 627 -836 631 -676
rect 652 -717 656 -677
rect 660 -717 664 -677
rect 850 -883 854 -843
rect 858 -883 862 -843
rect 902 -883 906 -843
rect 910 -883 914 -843
rect 954 -885 958 -845
rect 962 -885 966 -845
rect 980 -884 984 -843
rect 988 -884 992 -843
rect 997 -883 1001 -843
rect 1005 -883 1009 -843
rect 1019 -883 1023 -843
rect 1027 -883 1031 -843
rect 1131 -883 1135 -843
rect 1139 -883 1143 -843
rect 718 -1020 722 -980
rect 726 -1020 730 -980
rect 762 -986 766 -946
rect 770 -986 774 -946
rect 792 -986 796 -946
rect 800 -986 804 -946
rect 846 -988 850 -949
rect 854 -988 858 -949
rect 913 -982 917 -943
rect 921 -982 925 -943
rect -96 -1096 -56 -1092
rect -96 -1104 -56 -1100
rect -96 -1113 -55 -1109
rect -96 -1121 -55 -1117
rect -94 -1139 -54 -1135
rect -94 -1147 -54 -1143
rect 4 -1180 43 -1176
rect -96 -1191 -56 -1187
rect 4 -1188 43 -1184
rect -96 -1199 -56 -1195
rect -96 -1243 -56 -1239
rect -96 -1251 -56 -1247
rect 10 -1247 49 -1243
rect 10 -1255 49 -1251
rect -106 -1382 -102 -1342
rect -98 -1382 -94 -1342
rect -54 -1382 -50 -1342
rect -46 -1382 -42 -1342
rect -2 -1384 2 -1344
rect 6 -1384 10 -1344
rect 24 -1383 28 -1342
rect 32 -1383 36 -1342
rect 41 -1382 45 -1342
rect 49 -1382 53 -1342
rect 63 -1382 67 -1342
rect 71 -1382 75 -1342
rect 165 -1377 169 -1337
rect 173 -1377 177 -1337
rect 209 -1343 213 -1303
rect 217 -1343 221 -1303
rect 239 -1343 243 -1303
rect 247 -1343 251 -1303
rect 499 -1355 503 -1155
rect 507 -1355 511 -1155
rect 518 -1355 522 -1155
rect 526 -1355 530 -1155
rect 536 -1355 540 -1155
rect 544 -1355 548 -1155
rect 554 -1255 558 -1155
rect 562 -1255 566 -1155
rect -110 -1487 -106 -1448
rect -102 -1487 -98 -1448
rect -43 -1481 -39 -1442
rect -35 -1481 -31 -1442
rect 171 -1509 175 -1469
rect 179 -1509 183 -1469
rect 190 -1509 194 -1469
rect 198 -1509 202 -1469
rect 225 -1509 229 -1469
rect 233 -1509 237 -1469
rect 72 -1614 112 -1610
rect 72 -1622 112 -1618
rect 571 -1355 575 -1155
rect 579 -1355 583 -1155
rect 589 -1221 593 -1155
rect 597 -1221 601 -1155
rect 607 -1355 611 -1155
rect 615 -1355 619 -1155
rect 626 -1205 630 -1155
rect 634 -1205 638 -1155
rect 645 -1355 649 -1155
rect 653 -1355 657 -1155
rect 681 -1209 685 -1169
rect 689 -1209 693 -1169
rect 743 -1315 747 -1275
rect 751 -1315 755 -1275
rect 795 -1315 799 -1275
rect 803 -1315 807 -1275
rect 847 -1317 851 -1277
rect 855 -1317 859 -1277
rect 873 -1316 877 -1275
rect 881 -1316 885 -1275
rect 890 -1315 894 -1275
rect 898 -1315 902 -1275
rect 912 -1315 916 -1275
rect 920 -1315 924 -1275
rect 1024 -1315 1028 -1275
rect 1032 -1315 1036 -1275
rect 739 -1420 743 -1381
rect 747 -1420 751 -1381
rect 806 -1414 810 -1375
rect 814 -1414 818 -1375
rect 72 -1636 112 -1632
rect 72 -1644 112 -1640
rect 72 -1653 113 -1649
rect 72 -1661 113 -1657
rect 74 -1679 114 -1675
rect 74 -1687 114 -1683
rect 172 -1720 211 -1716
rect 72 -1731 112 -1727
rect 172 -1728 211 -1724
rect 72 -1739 112 -1735
rect 72 -1783 112 -1779
rect 72 -1791 112 -1787
rect 178 -1787 217 -1783
rect 178 -1795 217 -1791
<< polysilicon >>
rect 315 220 329 222
rect 349 220 352 222
rect 372 220 400 222
rect 439 220 442 222
rect 483 216 505 218
rect 545 216 548 218
rect 798 214 800 217
rect 850 214 852 217
rect 14 199 28 201
rect 48 199 51 201
rect 71 199 99 201
rect 138 199 141 201
rect 182 195 204 197
rect 244 195 247 197
rect 902 212 904 215
rect 928 214 930 217
rect 945 214 947 217
rect 967 214 969 217
rect 1058 214 1060 217
rect 364 172 461 174
rect 364 162 366 172
rect 459 166 461 172
rect 459 164 505 166
rect 545 164 548 166
rect 315 160 329 162
rect 349 160 366 162
rect 376 153 406 155
rect 445 153 448 155
rect 63 151 160 153
rect 63 141 65 151
rect 158 145 160 151
rect 798 152 800 174
rect 158 143 204 145
rect 244 143 247 145
rect 14 139 28 141
rect 48 139 65 141
rect 75 132 105 134
rect 144 132 147 134
rect 850 130 852 174
rect 842 128 852 130
rect 902 129 904 172
rect 364 120 460 122
rect 364 117 366 120
rect 317 115 330 117
rect 350 115 366 117
rect 458 114 460 120
rect 458 112 503 114
rect 543 112 546 114
rect 375 109 396 111
rect 416 109 419 111
rect 794 108 796 111
rect 63 99 159 101
rect 63 96 65 99
rect 16 94 29 96
rect 49 94 65 96
rect 157 93 159 99
rect 354 98 434 100
rect 157 91 202 93
rect 242 91 245 93
rect 74 88 95 90
rect 115 88 118 90
rect 354 88 356 98
rect 315 86 330 88
rect 350 86 356 88
rect 432 88 434 98
rect 377 86 397 88
rect 417 86 420 88
rect 432 86 504 88
rect 545 86 548 88
rect 53 77 133 79
rect -201 70 -199 73
rect -149 70 -147 73
rect -97 68 -95 71
rect -71 70 -69 73
rect -54 70 -52 73
rect -32 70 -30 73
rect -201 8 -199 30
rect -149 -14 -147 30
rect 53 67 55 77
rect 14 65 29 67
rect 49 65 55 67
rect 131 67 133 77
rect 393 69 397 71
rect 417 69 505 71
rect 545 69 548 71
rect 76 65 96 67
rect 116 65 119 67
rect 131 65 203 67
rect 244 65 247 67
rect 92 48 96 50
rect 116 48 204 50
rect 244 48 247 50
rect 394 47 397 49
rect 417 47 505 49
rect 545 47 548 49
rect 715 39 717 46
rect 745 39 747 42
rect 794 41 796 69
rect -157 -16 -147 -14
rect -97 -15 -95 28
rect -205 -36 -203 -33
rect -205 -103 -203 -75
rect -157 -109 -155 -16
rect -105 -17 -95 -15
rect -138 -30 -136 -27
rect -138 -99 -136 -69
rect -105 -109 -103 -17
rect -71 -41 -69 29
rect -83 -43 -69 -41
rect -94 -59 -92 -56
rect -94 -100 -92 -79
rect -157 -111 -143 -109
rect -105 -111 -98 -109
rect -205 -126 -203 -123
rect -145 -126 -143 -111
rect -100 -125 -98 -111
rect -83 -119 -81 -43
rect -71 -58 -69 -55
rect -54 -58 -52 30
rect -32 -58 -30 30
rect 93 26 96 28
rect 116 26 204 28
rect 244 26 247 28
rect 671 5 673 8
rect 189 -31 191 -24
rect 219 -31 221 -28
rect 145 -65 147 -62
rect -71 -98 -69 -78
rect -54 -82 -52 -78
rect -32 -81 -30 -78
rect 842 35 844 128
rect 894 127 904 129
rect 861 114 863 117
rect 861 45 863 75
rect 894 35 896 127
rect 928 103 930 173
rect 916 101 930 103
rect 905 85 907 88
rect 905 44 907 65
rect 842 33 856 35
rect 894 33 901 35
rect 794 18 796 21
rect 854 18 856 33
rect 899 19 901 33
rect 916 25 918 101
rect 928 86 930 89
rect 945 86 947 174
rect 967 86 969 174
rect 1058 86 1060 174
rect 928 46 930 66
rect 945 62 947 66
rect 967 63 969 66
rect 1058 63 1060 66
rect 916 23 930 25
rect 928 19 930 23
rect 715 -4 717 -1
rect 715 -24 717 -21
rect 745 -24 747 -1
rect 794 -16 796 -2
rect 854 -16 856 -2
rect 899 -14 901 -1
rect 928 -16 930 -1
rect 510 -40 512 -37
rect 527 -40 529 -37
rect 558 -40 560 -37
rect 189 -74 191 -71
rect 189 -94 191 -91
rect 219 -94 221 -71
rect -83 -121 -69 -119
rect -71 -125 -69 -121
rect 145 -128 147 -105
rect 189 -120 191 -113
rect 219 -117 221 -113
rect 600 -42 602 -39
rect 671 -58 673 -35
rect 715 -50 717 -43
rect 745 -47 747 -43
rect 671 -81 673 -77
rect 788 -82 790 -79
rect 840 -82 842 -79
rect -205 -160 -203 -146
rect -145 -160 -143 -146
rect -100 -158 -98 -145
rect -71 -160 -69 -145
rect 145 -151 147 -147
rect 151 -197 153 -194
rect 170 -197 172 -194
rect 205 -197 207 -194
rect -184 -217 -170 -215
rect -150 -217 -147 -215
rect -127 -217 -99 -215
rect -60 -217 -57 -215
rect -16 -221 6 -219
rect 46 -221 49 -219
rect 510 -211 512 -120
rect 527 -211 529 -120
rect -135 -265 -38 -263
rect -135 -275 -133 -265
rect -40 -271 -38 -265
rect 151 -269 153 -237
rect 170 -269 172 -237
rect 205 -262 207 -237
rect 558 -230 560 -120
rect 600 -227 602 -82
rect 892 -84 894 -81
rect 918 -82 920 -79
rect 935 -82 937 -79
rect 957 -82 959 -79
rect 1069 -82 1071 -79
rect 788 -144 790 -122
rect 840 -166 842 -122
rect 700 -173 702 -166
rect 832 -168 842 -166
rect 892 -167 894 -124
rect 730 -173 732 -170
rect 656 -207 658 -204
rect 784 -188 786 -185
rect 700 -216 702 -213
rect 700 -236 702 -233
rect 730 -236 732 -213
rect 510 -254 512 -251
rect 527 -254 529 -251
rect 558 -253 560 -250
rect 600 -252 602 -247
rect -40 -273 6 -271
rect 46 -273 49 -271
rect -184 -277 -170 -275
rect -150 -277 -133 -275
rect -123 -284 -93 -282
rect -54 -284 -51 -282
rect 656 -270 658 -247
rect 784 -255 786 -227
rect 700 -262 702 -255
rect 730 -259 732 -255
rect 832 -261 834 -168
rect 884 -169 894 -167
rect 851 -182 853 -179
rect 851 -251 853 -221
rect 884 -261 886 -169
rect 918 -193 920 -123
rect 906 -195 920 -193
rect 895 -211 897 -208
rect 895 -252 897 -231
rect 832 -263 846 -261
rect 884 -263 891 -261
rect 205 -286 207 -282
rect 784 -278 786 -275
rect 844 -278 846 -263
rect 889 -277 891 -263
rect 906 -271 908 -195
rect 918 -210 920 -207
rect 935 -210 937 -122
rect 957 -210 959 -122
rect 1069 -210 1071 -122
rect 918 -250 920 -230
rect 935 -234 937 -230
rect 957 -233 959 -230
rect 1069 -233 1071 -230
rect 906 -273 920 -271
rect 918 -277 920 -273
rect 656 -293 658 -289
rect 151 -313 153 -309
rect 170 -313 172 -309
rect 784 -312 786 -298
rect 844 -312 846 -298
rect 889 -310 891 -297
rect 918 -312 920 -297
rect -135 -317 -39 -315
rect -135 -320 -133 -317
rect -182 -322 -169 -320
rect -149 -322 -133 -320
rect -41 -323 -39 -317
rect -41 -325 4 -323
rect 44 -325 47 -323
rect -124 -328 -103 -326
rect -83 -328 -80 -326
rect -145 -339 -65 -337
rect -145 -349 -143 -339
rect -184 -351 -169 -349
rect -149 -351 -143 -349
rect -67 -349 -65 -339
rect 211 -345 213 -338
rect 241 -345 243 -342
rect -122 -351 -102 -349
rect -82 -351 -79 -349
rect -67 -351 5 -349
rect 46 -351 49 -349
rect -106 -368 -102 -366
rect -82 -368 6 -366
rect 46 -368 49 -366
rect 167 -379 169 -376
rect -105 -390 -102 -388
rect -82 -390 6 -388
rect 46 -390 49 -388
rect 515 -371 517 -368
rect 527 -371 529 -368
rect 211 -388 213 -385
rect 211 -408 213 -405
rect 241 -408 243 -385
rect 167 -442 169 -419
rect 211 -434 213 -427
rect 241 -431 243 -427
rect -119 -453 -117 -450
rect -67 -453 -65 -450
rect -15 -455 -13 -452
rect 11 -453 13 -450
rect 28 -453 30 -450
rect 50 -453 52 -450
rect -119 -515 -117 -493
rect -67 -537 -65 -493
rect 167 -465 169 -461
rect 546 -372 548 -368
rect 564 -372 566 -369
rect 583 -372 585 -369
rect -75 -539 -65 -537
rect -15 -538 -13 -495
rect -123 -559 -121 -556
rect -123 -626 -121 -598
rect -75 -632 -73 -539
rect -23 -540 -13 -538
rect -56 -553 -54 -550
rect -56 -622 -54 -592
rect -23 -632 -21 -540
rect 11 -564 13 -494
rect -1 -566 13 -564
rect -12 -582 -10 -579
rect -12 -623 -10 -602
rect -75 -634 -61 -632
rect -23 -634 -16 -632
rect -123 -649 -121 -646
rect -63 -649 -61 -634
rect -18 -648 -16 -634
rect -1 -642 1 -566
rect 11 -581 13 -578
rect 28 -581 30 -493
rect 50 -581 52 -493
rect 173 -511 175 -508
rect 192 -511 194 -508
rect 227 -511 229 -508
rect 173 -583 175 -551
rect 192 -583 194 -551
rect 227 -576 229 -551
rect 515 -570 517 -491
rect 527 -570 529 -491
rect 668 -383 670 -368
rect 862 -415 864 -412
rect 914 -415 916 -412
rect 668 -459 670 -423
rect 776 -429 778 -422
rect 806 -429 808 -426
rect 732 -463 734 -460
rect 668 -482 670 -479
rect 546 -570 548 -492
rect 564 -570 566 -492
rect 583 -570 585 -492
rect 966 -417 968 -414
rect 992 -415 994 -412
rect 1009 -415 1011 -412
rect 1031 -415 1033 -412
rect 1136 -415 1138 -412
rect 776 -472 778 -469
rect 776 -492 778 -489
rect 806 -492 808 -469
rect 862 -477 864 -455
rect 732 -526 734 -503
rect 914 -499 916 -455
rect 906 -501 916 -499
rect 966 -500 968 -457
rect 776 -518 778 -511
rect 806 -515 808 -511
rect 858 -521 860 -518
rect 732 -549 734 -545
rect 11 -621 13 -601
rect 28 -605 30 -601
rect 50 -604 52 -601
rect 227 -600 229 -596
rect 173 -627 175 -623
rect 192 -627 194 -623
rect 546 -604 548 -600
rect 858 -588 860 -560
rect 583 -594 585 -590
rect 906 -594 908 -501
rect 958 -502 968 -500
rect 925 -515 927 -512
rect 925 -584 927 -554
rect 958 -594 960 -502
rect 992 -526 994 -456
rect 980 -528 994 -526
rect 969 -544 971 -541
rect 969 -585 971 -564
rect 906 -596 920 -594
rect 958 -596 965 -594
rect 858 -611 860 -608
rect 918 -611 920 -596
rect 963 -610 965 -596
rect 980 -604 982 -528
rect 992 -543 994 -540
rect 1009 -543 1011 -455
rect 1031 -543 1033 -455
rect 1136 -543 1138 -455
rect 992 -583 994 -563
rect 1009 -567 1011 -563
rect 1031 -566 1033 -563
rect 1136 -566 1138 -563
rect 980 -606 994 -604
rect 992 -610 994 -606
rect 515 -633 517 -630
rect 527 -633 529 -630
rect 564 -633 566 -630
rect -1 -644 13 -642
rect 11 -648 13 -644
rect 858 -645 860 -631
rect 918 -645 920 -631
rect 963 -643 965 -630
rect 992 -645 994 -630
rect -123 -683 -121 -669
rect -63 -683 -61 -669
rect -18 -681 -16 -668
rect 11 -683 13 -668
rect 514 -678 516 -675
rect 532 -678 534 -675
rect 550 -678 552 -675
rect 568 -678 570 -675
rect 587 -677 589 -674
rect 606 -677 608 -674
rect 624 -676 626 -673
rect -99 -732 -97 -729
rect -47 -732 -45 -729
rect 5 -734 7 -731
rect 31 -732 33 -729
rect 48 -732 50 -729
rect 70 -732 72 -729
rect -99 -794 -97 -772
rect -47 -816 -45 -772
rect -55 -818 -45 -816
rect 5 -817 7 -774
rect -103 -838 -101 -835
rect -103 -905 -101 -877
rect -55 -911 -53 -818
rect -3 -819 7 -817
rect -36 -832 -34 -829
rect -36 -901 -34 -871
rect -3 -911 -1 -819
rect 31 -843 33 -773
rect 19 -845 33 -843
rect 8 -861 10 -858
rect 8 -902 10 -881
rect -55 -913 -41 -911
rect -3 -913 4 -911
rect -103 -928 -101 -925
rect -43 -928 -41 -913
rect 2 -927 4 -913
rect 19 -921 21 -845
rect 31 -860 33 -857
rect 48 -860 50 -772
rect 70 -860 72 -772
rect 211 -774 213 -767
rect 241 -774 243 -771
rect 167 -808 169 -805
rect 211 -817 213 -814
rect 211 -837 213 -834
rect 241 -837 243 -814
rect 167 -871 169 -848
rect 211 -863 213 -856
rect 241 -860 243 -856
rect 31 -900 33 -880
rect 48 -884 50 -880
rect 70 -883 72 -880
rect 167 -894 169 -890
rect 19 -923 33 -921
rect 31 -927 33 -923
rect 173 -940 175 -937
rect 192 -940 194 -937
rect 227 -940 229 -937
rect -103 -962 -101 -948
rect -43 -962 -41 -948
rect 2 -960 4 -947
rect 31 -962 33 -947
rect 173 -1012 175 -980
rect 192 -1012 194 -980
rect 227 -1005 229 -980
rect 514 -1008 516 -838
rect 227 -1029 229 -1025
rect 173 -1056 175 -1052
rect 192 -1056 194 -1052
rect -99 -1077 -96 -1075
rect -56 -1077 32 -1075
rect 52 -1077 55 -1075
rect 532 -1009 534 -838
rect 514 -1091 516 -1088
rect 550 -1048 552 -838
rect 568 -1009 570 -758
rect 532 -1092 534 -1089
rect 550 -1092 552 -1088
rect 587 -1062 589 -837
rect 606 -1008 608 -731
rect 657 -677 659 -674
rect 624 -1068 626 -836
rect 657 -1068 659 -717
rect 855 -843 857 -840
rect 907 -843 909 -840
rect 959 -845 961 -842
rect 985 -843 987 -840
rect 1002 -843 1004 -840
rect 1024 -843 1026 -840
rect 1136 -843 1138 -840
rect 855 -905 857 -883
rect 907 -927 909 -883
rect 899 -929 909 -927
rect 959 -928 961 -885
rect 767 -946 769 -939
rect 797 -946 799 -943
rect 723 -980 725 -977
rect 851 -949 853 -946
rect 767 -989 769 -986
rect 767 -1009 769 -1006
rect 797 -1009 799 -986
rect 723 -1043 725 -1020
rect 851 -1016 853 -988
rect 899 -1022 901 -929
rect 951 -930 961 -928
rect 918 -943 920 -940
rect 918 -1012 920 -982
rect 951 -1022 953 -930
rect 985 -954 987 -884
rect 973 -956 987 -954
rect 962 -972 964 -969
rect 962 -1013 964 -992
rect 899 -1024 913 -1022
rect 951 -1024 958 -1022
rect 767 -1035 769 -1028
rect 797 -1032 799 -1028
rect 851 -1039 853 -1036
rect 911 -1039 913 -1024
rect 956 -1038 958 -1024
rect 973 -1032 975 -956
rect 985 -971 987 -968
rect 1002 -971 1004 -883
rect 1024 -971 1026 -883
rect 1136 -971 1138 -883
rect 985 -1011 987 -991
rect 1002 -995 1004 -991
rect 1024 -994 1026 -991
rect 1136 -994 1138 -991
rect 973 -1034 987 -1032
rect 985 -1038 987 -1034
rect 723 -1066 725 -1062
rect 851 -1073 853 -1059
rect 911 -1073 913 -1059
rect 956 -1071 958 -1058
rect 985 -1073 987 -1058
rect 568 -1092 570 -1089
rect 587 -1091 589 -1088
rect 606 -1092 608 -1088
rect 624 -1092 626 -1088
rect 657 -1091 659 -1088
rect -99 -1099 -96 -1097
rect -56 -1099 32 -1097
rect 52 -1099 56 -1097
rect -99 -1116 -96 -1114
rect -55 -1116 17 -1114
rect 29 -1116 32 -1114
rect 52 -1116 72 -1114
rect 15 -1126 17 -1116
rect 93 -1116 99 -1114
rect 119 -1116 134 -1114
rect 93 -1126 95 -1116
rect 15 -1128 95 -1126
rect 30 -1139 33 -1137
rect 53 -1139 74 -1137
rect -97 -1142 -94 -1140
rect -54 -1142 -9 -1140
rect -11 -1148 -9 -1142
rect 83 -1145 99 -1143
rect 119 -1145 132 -1143
rect 83 -1148 85 -1145
rect -11 -1150 85 -1148
rect 504 -1155 506 -1152
rect 523 -1155 525 -1151
rect 541 -1155 543 -1151
rect 559 -1155 561 -1151
rect 576 -1155 578 -1152
rect 594 -1155 596 -1151
rect 612 -1155 614 -1152
rect 631 -1155 633 -1152
rect 650 -1155 652 -1152
rect 1 -1183 4 -1181
rect 43 -1183 73 -1181
rect 83 -1190 100 -1188
rect 120 -1190 134 -1188
rect -99 -1194 -96 -1192
rect -56 -1194 -10 -1192
rect -12 -1200 -10 -1194
rect 83 -1200 85 -1190
rect -12 -1202 85 -1200
rect -99 -1246 -96 -1244
rect -56 -1246 -34 -1244
rect 7 -1250 10 -1248
rect 49 -1250 77 -1248
rect 97 -1250 100 -1248
rect 120 -1250 134 -1248
rect 214 -1303 216 -1296
rect 244 -1303 246 -1300
rect 170 -1337 172 -1334
rect -101 -1342 -99 -1339
rect -49 -1342 -47 -1339
rect 3 -1344 5 -1341
rect 29 -1342 31 -1339
rect 46 -1342 48 -1339
rect 68 -1342 70 -1339
rect -101 -1404 -99 -1382
rect -49 -1426 -47 -1382
rect 214 -1346 216 -1343
rect 214 -1366 216 -1363
rect 244 -1366 246 -1343
rect -57 -1428 -47 -1426
rect 3 -1427 5 -1384
rect -105 -1448 -103 -1445
rect -105 -1515 -103 -1487
rect -57 -1521 -55 -1428
rect -5 -1429 5 -1427
rect -38 -1442 -36 -1439
rect -38 -1511 -36 -1481
rect -5 -1521 -3 -1429
rect 29 -1453 31 -1383
rect 17 -1455 31 -1453
rect 6 -1471 8 -1468
rect 6 -1512 8 -1491
rect -57 -1523 -43 -1521
rect -5 -1523 2 -1521
rect -105 -1538 -103 -1535
rect -45 -1538 -43 -1523
rect 0 -1537 2 -1523
rect 17 -1531 19 -1455
rect 29 -1470 31 -1467
rect 46 -1470 48 -1382
rect 68 -1470 70 -1382
rect 170 -1400 172 -1377
rect 214 -1392 216 -1385
rect 244 -1389 246 -1385
rect 170 -1423 172 -1419
rect 176 -1469 178 -1466
rect 195 -1469 197 -1466
rect 230 -1469 232 -1466
rect 29 -1510 31 -1490
rect 46 -1494 48 -1490
rect 68 -1493 70 -1490
rect 17 -1533 31 -1531
rect 29 -1537 31 -1533
rect 176 -1541 178 -1509
rect 195 -1541 197 -1509
rect 230 -1534 232 -1509
rect 504 -1532 506 -1355
rect 523 -1532 525 -1355
rect -105 -1572 -103 -1558
rect -45 -1572 -43 -1558
rect 0 -1570 2 -1557
rect 29 -1572 31 -1557
rect 230 -1558 232 -1554
rect 176 -1585 178 -1581
rect 195 -1585 197 -1581
rect 69 -1617 72 -1615
rect 112 -1617 200 -1615
rect 220 -1617 223 -1615
rect 541 -1582 543 -1355
rect 559 -1532 561 -1255
rect 576 -1599 578 -1355
rect 594 -1532 596 -1221
rect 612 -1607 614 -1355
rect 631 -1532 633 -1205
rect 686 -1169 688 -1166
rect 650 -1612 652 -1355
rect 686 -1612 688 -1209
rect 748 -1275 750 -1272
rect 800 -1275 802 -1272
rect 852 -1277 854 -1274
rect 878 -1275 880 -1272
rect 895 -1275 897 -1272
rect 917 -1275 919 -1272
rect 1029 -1275 1031 -1272
rect 748 -1337 750 -1315
rect 800 -1359 802 -1315
rect 792 -1361 802 -1359
rect 852 -1360 854 -1317
rect 744 -1381 746 -1378
rect 744 -1448 746 -1420
rect 792 -1454 794 -1361
rect 844 -1362 854 -1360
rect 811 -1375 813 -1372
rect 811 -1444 813 -1414
rect 844 -1454 846 -1362
rect 878 -1386 880 -1316
rect 866 -1388 880 -1386
rect 855 -1404 857 -1401
rect 855 -1445 857 -1424
rect 792 -1456 806 -1454
rect 844 -1456 851 -1454
rect 744 -1471 746 -1468
rect 804 -1471 806 -1456
rect 849 -1470 851 -1456
rect 866 -1464 868 -1388
rect 878 -1403 880 -1400
rect 895 -1403 897 -1315
rect 917 -1403 919 -1315
rect 1029 -1403 1031 -1315
rect 878 -1443 880 -1423
rect 895 -1427 897 -1423
rect 917 -1426 919 -1423
rect 1029 -1426 1031 -1423
rect 866 -1466 880 -1464
rect 878 -1470 880 -1466
rect 744 -1505 746 -1491
rect 804 -1505 806 -1491
rect 849 -1503 851 -1490
rect 878 -1505 880 -1490
rect 504 -1635 506 -1632
rect 523 -1635 525 -1632
rect 541 -1635 543 -1632
rect 559 -1635 561 -1632
rect 576 -1635 578 -1632
rect 594 -1635 596 -1632
rect 612 -1635 614 -1632
rect 631 -1635 633 -1632
rect 650 -1635 652 -1632
rect 686 -1635 688 -1632
rect 69 -1639 72 -1637
rect 112 -1639 200 -1637
rect 220 -1639 224 -1637
rect 69 -1656 72 -1654
rect 113 -1656 185 -1654
rect 197 -1656 200 -1654
rect 220 -1656 240 -1654
rect 183 -1666 185 -1656
rect 261 -1656 267 -1654
rect 287 -1656 302 -1654
rect 261 -1666 263 -1656
rect 183 -1668 263 -1666
rect 198 -1679 201 -1677
rect 221 -1679 242 -1677
rect 71 -1682 74 -1680
rect 114 -1682 159 -1680
rect 157 -1688 159 -1682
rect 251 -1685 267 -1683
rect 287 -1685 300 -1683
rect 251 -1688 253 -1685
rect 157 -1690 253 -1688
rect 169 -1723 172 -1721
rect 211 -1723 241 -1721
rect 251 -1730 268 -1728
rect 288 -1730 302 -1728
rect 69 -1734 72 -1732
rect 112 -1734 158 -1732
rect 156 -1740 158 -1734
rect 251 -1740 253 -1730
rect 156 -1742 253 -1740
rect 69 -1786 72 -1784
rect 112 -1786 134 -1784
rect 175 -1790 178 -1788
rect 217 -1790 245 -1788
rect 265 -1790 268 -1788
rect 288 -1790 302 -1788
<< polycontact >>
rect 316 222 320 226
rect 372 222 376 226
rect 483 218 487 222
rect 15 201 19 205
rect 71 201 75 205
rect 182 197 186 201
rect 485 166 489 170
rect 376 155 380 159
rect 794 152 798 156
rect 846 154 850 158
rect 184 145 188 149
rect 75 134 79 138
rect 898 139 902 143
rect 924 139 928 143
rect 375 111 379 115
rect 470 114 474 118
rect 74 90 78 94
rect 169 93 173 97
rect 377 88 381 92
rect 470 88 474 92
rect -205 8 -201 12
rect -153 10 -149 14
rect 76 67 80 71
rect 169 67 173 71
rect 470 71 474 75
rect 169 50 173 54
rect 470 49 474 53
rect 711 42 715 46
rect 790 41 794 45
rect -101 -5 -97 -1
rect -75 -5 -71 -1
rect -209 -103 -205 -99
rect -142 -99 -138 -95
rect -58 -5 -54 -1
rect -98 -100 -94 -96
rect -36 -5 -32 -1
rect 169 28 173 32
rect 185 -28 189 -24
rect -75 -98 -71 -94
rect 857 45 861 49
rect 941 139 945 143
rect 901 44 905 48
rect 963 139 967 143
rect 1054 139 1058 143
rect 924 46 928 50
rect 741 -16 745 -12
rect 790 -15 794 -11
rect 215 -86 219 -82
rect 141 -120 145 -116
rect 185 -120 189 -116
rect 667 -50 671 -46
rect 711 -50 715 -46
rect -209 -159 -205 -155
rect 506 -137 510 -133
rect -183 -215 -179 -211
rect -127 -215 -123 -211
rect -16 -219 -12 -215
rect 523 -175 527 -171
rect 554 -208 558 -204
rect 147 -248 151 -244
rect -14 -271 -10 -267
rect 166 -258 170 -254
rect 201 -248 205 -244
rect 596 -172 600 -167
rect 784 -144 788 -140
rect 836 -142 840 -138
rect 888 -157 892 -153
rect 696 -170 700 -166
rect 914 -157 918 -153
rect 726 -228 730 -224
rect 652 -262 656 -258
rect -123 -282 -119 -278
rect 780 -255 784 -251
rect 696 -262 700 -258
rect 847 -251 851 -247
rect 931 -157 935 -153
rect 891 -252 895 -248
rect 953 -157 957 -153
rect 1065 -157 1069 -153
rect 914 -250 918 -246
rect 780 -311 784 -307
rect -124 -326 -120 -322
rect -29 -323 -25 -319
rect -122 -349 -118 -345
rect 207 -342 211 -338
rect -29 -349 -25 -345
rect -29 -366 -25 -362
rect -29 -388 -25 -384
rect 237 -400 241 -396
rect 163 -434 167 -430
rect 207 -434 211 -430
rect -123 -515 -119 -511
rect -71 -513 -67 -509
rect -19 -528 -15 -524
rect 7 -528 11 -524
rect -127 -626 -123 -622
rect -60 -622 -56 -618
rect 24 -528 28 -524
rect -16 -623 -12 -619
rect 46 -528 50 -524
rect 511 -507 515 -503
rect 169 -562 173 -558
rect 188 -572 192 -568
rect 223 -562 227 -558
rect 523 -520 527 -516
rect 660 -450 668 -444
rect 772 -426 776 -422
rect 542 -534 546 -530
rect 560 -548 564 -544
rect 579 -559 583 -555
rect 802 -484 806 -480
rect 858 -477 862 -473
rect 910 -475 914 -471
rect 728 -518 732 -514
rect 962 -490 966 -486
rect 988 -490 992 -486
rect 772 -518 776 -514
rect 7 -621 11 -617
rect 854 -588 858 -584
rect 921 -584 925 -580
rect 1005 -490 1009 -486
rect 965 -585 969 -581
rect 1027 -490 1031 -486
rect 1132 -490 1136 -486
rect 988 -583 992 -579
rect 854 -644 858 -640
rect -127 -682 -123 -678
rect -103 -794 -99 -790
rect -51 -792 -47 -788
rect 207 -771 211 -767
rect 1 -807 5 -803
rect 27 -807 31 -803
rect -107 -905 -103 -901
rect -40 -901 -36 -897
rect 44 -807 48 -803
rect 4 -902 8 -898
rect 66 -807 70 -803
rect 237 -829 241 -825
rect 163 -863 167 -859
rect 509 -855 514 -848
rect 207 -863 211 -859
rect 27 -900 31 -896
rect -107 -961 -103 -957
rect 169 -991 173 -987
rect 188 -1001 192 -997
rect 223 -991 227 -987
rect 527 -874 532 -867
rect -25 -1081 -21 -1077
rect 545 -892 550 -885
rect 563 -913 568 -906
rect 582 -935 587 -928
rect 601 -962 606 -955
rect 619 -991 624 -984
rect 653 -966 657 -962
rect 851 -905 855 -901
rect 903 -903 907 -899
rect 955 -918 959 -914
rect 981 -918 985 -914
rect 763 -943 767 -939
rect 793 -1001 797 -997
rect 719 -1035 723 -1031
rect 847 -1016 851 -1012
rect 914 -1012 918 -1008
rect 998 -918 1002 -914
rect 958 -1013 962 -1009
rect 763 -1035 767 -1031
rect 1020 -918 1024 -914
rect 1132 -918 1136 -914
rect 981 -1011 985 -1007
rect 847 -1072 851 -1068
rect -25 -1103 -21 -1099
rect -25 -1120 -21 -1116
rect 68 -1120 72 -1116
rect -25 -1146 -21 -1142
rect 70 -1143 74 -1139
rect 69 -1187 73 -1183
rect -40 -1198 -36 -1194
rect -38 -1250 -34 -1246
rect 73 -1254 77 -1250
rect 129 -1254 133 -1250
rect 210 -1300 214 -1296
rect -105 -1404 -101 -1400
rect -53 -1402 -49 -1398
rect 240 -1358 244 -1354
rect -1 -1417 3 -1413
rect 25 -1417 29 -1413
rect -109 -1515 -105 -1511
rect -42 -1511 -38 -1507
rect 42 -1417 46 -1413
rect 2 -1512 6 -1508
rect 64 -1417 68 -1413
rect 166 -1392 170 -1388
rect 210 -1392 214 -1388
rect 499 -1399 504 -1394
rect 25 -1510 29 -1506
rect 172 -1520 176 -1516
rect 191 -1530 195 -1526
rect 226 -1520 230 -1516
rect 518 -1413 523 -1408
rect 536 -1430 541 -1425
rect -109 -1571 -105 -1567
rect 143 -1621 147 -1617
rect 554 -1444 559 -1439
rect 571 -1460 576 -1455
rect 589 -1473 594 -1468
rect 607 -1490 612 -1485
rect 626 -1504 631 -1499
rect 645 -1520 650 -1515
rect 681 -1409 686 -1403
rect 744 -1337 748 -1333
rect 796 -1335 800 -1331
rect 848 -1350 852 -1346
rect 874 -1350 878 -1346
rect 740 -1448 744 -1444
rect 807 -1444 811 -1440
rect 891 -1350 895 -1346
rect 851 -1445 855 -1441
rect 913 -1350 917 -1346
rect 1025 -1350 1029 -1346
rect 874 -1443 878 -1439
rect 740 -1504 744 -1500
rect 143 -1643 147 -1639
rect 143 -1660 147 -1656
rect 236 -1660 240 -1656
rect 143 -1686 147 -1682
rect 238 -1683 242 -1679
rect 237 -1727 241 -1723
rect 128 -1738 132 -1734
rect 130 -1790 134 -1786
rect 241 -1794 245 -1790
rect 297 -1794 301 -1790
<< polypplus >>
rect 564 -492 566 -432
<< metal1 >>
rect 387 250 392 251
rect 416 250 420 259
rect 316 245 487 250
rect 15 224 186 229
rect 1 198 11 207
rect 15 205 19 224
rect 48 202 57 206
rect 53 198 57 202
rect 71 205 75 212
rect 138 202 170 206
rect 1 194 28 198
rect 53 194 99 198
rect 166 194 170 202
rect 182 201 186 224
rect 302 219 312 228
rect 316 226 320 245
rect 349 223 358 227
rect 354 219 358 223
rect 372 226 376 233
rect 439 223 471 227
rect 251 202 269 217
rect 244 198 269 202
rect 1 138 11 194
rect 71 159 75 194
rect 166 190 204 194
rect 71 155 188 159
rect 184 149 188 155
rect 251 150 269 198
rect 48 142 59 146
rect 244 146 269 150
rect 1 134 28 138
rect -221 77 -14 95
rect 1 93 11 134
rect 55 131 59 142
rect 75 138 79 143
rect 171 139 204 142
rect 144 138 204 139
rect 144 135 177 138
rect 55 127 105 131
rect 75 109 79 127
rect 75 105 173 109
rect 49 97 58 101
rect 169 97 173 105
rect 251 98 269 146
rect 1 89 29 93
rect -206 70 -202 77
rect -154 70 -150 77
rect -233 8 -205 12
rect -233 -155 -228 8
rect -198 -4 -194 30
rect -210 -8 -194 -4
rect -163 10 -153 14
rect -210 -36 -206 -8
rect -202 -99 -198 -75
rect -163 -99 -159 10
rect -146 3 -142 30
rect -102 68 -98 77
rect -76 70 -72 77
rect -59 70 -55 77
rect -37 70 -33 77
rect -146 -3 -139 3
rect -94 -1 -90 28
rect -68 -1 -64 29
rect -51 -1 -47 30
rect -29 -1 -25 30
rect 1 64 11 89
rect 54 87 58 97
rect 74 94 78 97
rect 115 91 151 95
rect 242 94 269 98
rect 147 90 151 91
rect 54 83 95 87
rect 147 86 202 90
rect 49 68 62 72
rect 58 64 62 68
rect 76 71 80 74
rect 116 68 127 72
rect 123 64 127 68
rect 169 71 173 86
rect 251 72 269 94
rect 244 68 269 72
rect 1 60 29 64
rect 58 60 96 64
rect 123 60 203 64
rect 1 47 11 60
rect 116 51 129 55
rect 125 47 129 51
rect 169 54 173 60
rect 251 55 269 68
rect 244 51 269 55
rect 1 43 96 47
rect 125 43 204 47
rect 1 25 11 43
rect 116 29 127 33
rect 1 21 96 25
rect 123 21 127 29
rect 169 32 173 43
rect 251 33 269 51
rect 244 29 269 33
rect 167 21 204 25
rect 1 3 11 21
rect 123 17 173 21
rect -143 -30 -139 -3
rect -113 -5 -101 -1
rect -94 -5 -75 -1
rect -68 -5 -58 -1
rect -51 -5 -36 -1
rect -135 -95 -131 -69
rect -113 -95 -109 -5
rect -94 -23 -90 -5
rect -99 -27 -90 -23
rect -99 -59 -95 -27
rect -68 -47 -64 -5
rect -51 -45 -47 -5
rect -29 -7 -21 -1
rect -76 -51 -64 -47
rect -59 -49 -47 -45
rect -25 -47 -21 -7
rect 169 -16 173 17
rect 251 10 269 29
rect 302 215 329 219
rect 354 215 400 219
rect 467 215 471 223
rect 483 222 487 245
rect 552 223 570 238
rect 545 219 570 223
rect 778 221 985 239
rect 1046 221 1076 239
rect 302 159 312 215
rect 372 180 376 215
rect 467 211 505 215
rect 372 176 489 180
rect 485 170 489 176
rect 552 171 570 219
rect 793 214 797 221
rect 845 214 849 221
rect 349 163 360 167
rect 545 167 570 171
rect 302 155 329 159
rect 302 114 312 155
rect 356 152 360 163
rect 376 159 380 164
rect 472 160 505 163
rect 445 159 505 160
rect 445 156 478 159
rect 356 148 406 152
rect 376 130 380 148
rect 376 126 474 130
rect 350 118 359 122
rect 470 118 474 126
rect 552 119 570 167
rect 302 110 330 114
rect 302 85 312 110
rect 355 108 359 118
rect 375 115 379 118
rect 416 112 452 116
rect 543 115 570 119
rect 448 111 452 112
rect 355 104 396 108
rect 448 107 503 111
rect 350 89 363 93
rect 359 85 363 89
rect 377 92 381 95
rect 417 89 428 93
rect 424 85 428 89
rect 470 92 474 107
rect 552 93 570 115
rect 545 89 570 93
rect 302 81 330 85
rect 359 81 397 85
rect 424 81 504 85
rect 302 68 312 81
rect 417 72 430 76
rect 426 68 430 72
rect 470 75 474 81
rect 552 76 570 89
rect 545 72 570 76
rect 302 64 397 68
rect 426 64 505 68
rect 302 46 312 64
rect 417 50 428 54
rect 302 42 397 46
rect 424 42 428 50
rect 470 53 474 64
rect 552 54 570 72
rect 766 152 794 156
rect 545 50 570 54
rect 468 42 505 46
rect 302 24 312 42
rect 424 38 474 42
rect 470 24 474 38
rect 552 31 570 50
rect 691 49 744 54
rect 691 46 696 49
rect 652 42 711 46
rect 165 -21 218 -16
rect 165 -24 170 -21
rect 126 -28 185 -24
rect -76 -58 -72 -51
rect -59 -58 -55 -49
rect -37 -51 83 -47
rect -37 -58 -33 -51
rect -147 -99 -142 -95
rect -135 -99 -109 -95
rect -216 -103 -209 -99
rect -202 -103 -159 -99
rect -202 -117 -198 -103
rect -135 -115 -131 -99
rect -101 -100 -98 -96
rect -210 -121 -198 -117
rect -150 -119 -131 -115
rect -91 -116 -87 -79
rect -78 -98 -75 -94
rect -68 -112 -64 -78
rect -210 -126 -206 -121
rect -150 -126 -146 -119
rect -105 -120 -87 -116
rect -76 -116 -64 -112
rect -105 -125 -101 -120
rect -76 -125 -72 -116
rect -233 -159 -209 -155
rect -202 -163 -198 -146
rect -142 -163 -138 -146
rect -97 -163 -93 -145
rect -68 -163 -64 -145
rect -51 -163 -47 -78
rect -29 -163 -25 -78
rect 126 -116 131 -28
rect 214 -31 218 -21
rect 137 -60 154 -56
rect 140 -65 144 -60
rect 165 -82 170 -51
rect 184 -82 188 -71
rect 492 -33 614 -29
rect 192 -72 196 -71
rect 222 -81 226 -71
rect 505 -40 509 -33
rect 530 -40 534 -33
rect 165 -86 215 -82
rect 222 -86 231 -81
rect 236 -86 403 -81
rect 148 -116 152 -105
rect 184 -94 188 -86
rect 222 -94 226 -86
rect 104 -120 141 -116
rect 148 -120 185 -116
rect -211 -173 -7 -163
rect -183 -192 -12 -187
rect -197 -218 -187 -209
rect -183 -211 -179 -192
rect -150 -214 -141 -210
rect -145 -218 -141 -214
rect -127 -211 -123 -204
rect -60 -214 -28 -210
rect -197 -222 -170 -218
rect -145 -222 -99 -218
rect -32 -222 -28 -214
rect -16 -215 -12 -192
rect 53 -214 71 -199
rect 46 -218 71 -214
rect -197 -278 -187 -222
rect -127 -257 -123 -222
rect -32 -226 6 -222
rect -127 -261 -10 -257
rect -14 -267 -10 -261
rect 53 -266 71 -218
rect 104 -254 107 -120
rect 148 -128 152 -120
rect 172 -123 176 -120
rect 214 -123 218 -113
rect 172 -128 218 -123
rect 140 -153 144 -147
rect 135 -157 154 -153
rect 406 -171 410 -86
rect 517 -45 522 -40
rect 522 -123 526 -120
rect 553 -123 557 -120
rect 522 -128 557 -123
rect 595 -42 599 -33
rect 621 -46 624 -15
rect 652 -46 657 42
rect 740 39 744 49
rect 663 10 680 14
rect 666 5 670 10
rect 691 -12 696 19
rect 710 -12 714 -1
rect 718 -2 722 -1
rect 748 -11 752 -1
rect 766 -11 771 152
rect 801 140 805 174
rect 789 136 805 140
rect 836 154 846 158
rect 789 108 793 136
rect 797 45 801 69
rect 836 45 840 154
rect 853 147 857 174
rect 897 212 901 221
rect 923 214 927 221
rect 940 214 944 221
rect 962 214 966 221
rect 1053 214 1057 221
rect 853 141 860 147
rect 905 143 909 172
rect 931 143 935 173
rect 948 143 952 174
rect 970 143 974 174
rect 1061 143 1065 174
rect 856 114 860 141
rect 886 139 898 143
rect 905 139 924 143
rect 931 139 941 143
rect 948 139 963 143
rect 970 139 1054 143
rect 1061 139 1082 143
rect 864 49 868 75
rect 886 49 890 139
rect 905 121 909 139
rect 900 117 909 121
rect 900 85 904 117
rect 931 97 935 139
rect 948 99 952 139
rect 970 137 978 139
rect 1061 137 1069 139
rect 923 93 935 97
rect 940 95 952 99
rect 974 97 978 137
rect 1065 97 1069 137
rect 923 86 927 93
rect 940 86 944 95
rect 962 93 978 97
rect 1053 93 1069 97
rect 962 86 966 93
rect 1053 86 1057 93
rect 852 45 857 49
rect 864 45 890 49
rect 783 41 790 45
rect 797 41 840 45
rect 797 27 801 41
rect 864 29 868 45
rect 898 44 901 48
rect 789 23 801 27
rect 849 25 868 29
rect 908 28 912 65
rect 921 46 924 50
rect 931 32 935 66
rect 789 18 793 23
rect 849 18 853 25
rect 894 24 912 28
rect 923 28 935 32
rect 894 19 898 24
rect 923 19 927 28
rect 691 -16 741 -12
rect 748 -16 757 -11
rect 762 -15 790 -11
rect 762 -16 768 -15
rect 674 -46 678 -35
rect 710 -24 714 -16
rect 748 -24 752 -16
rect 797 -19 801 -2
rect 857 -19 861 -2
rect 902 -19 906 -1
rect 931 -19 935 -1
rect 948 -19 952 66
rect 970 -19 974 66
rect 1061 -19 1065 66
rect 788 -29 992 -19
rect 1046 -29 1082 -19
rect 621 -50 667 -46
rect 674 -50 711 -46
rect 674 -58 678 -50
rect 698 -53 702 -50
rect 740 -53 744 -43
rect 698 -58 744 -53
rect 768 -75 975 -57
rect 1057 -75 1087 -57
rect 666 -82 670 -77
rect 783 -82 787 -75
rect 835 -82 839 -75
rect 475 -137 506 -133
rect 561 -167 565 -120
rect 603 -131 607 -82
rect 661 -85 680 -82
rect 603 -135 634 -131
rect 406 -175 441 -171
rect 448 -175 523 -171
rect 561 -172 596 -167
rect 140 -190 219 -185
rect 146 -197 150 -190
rect 165 -197 169 -190
rect 200 -197 204 -190
rect 154 -244 158 -237
rect 173 -244 177 -237
rect 208 -244 212 -237
rect 477 -208 554 -204
rect 133 -248 147 -244
rect 159 -248 201 -244
rect 208 -248 406 -244
rect 208 -254 212 -248
rect 477 -244 482 -208
rect 412 -248 482 -244
rect 104 -258 166 -254
rect 200 -258 212 -254
rect 517 -216 522 -211
rect 561 -221 565 -172
rect 553 -225 565 -221
rect 553 -230 557 -225
rect 603 -227 607 -135
rect 629 -187 634 -135
rect 756 -144 784 -140
rect 676 -163 729 -158
rect 676 -166 681 -163
rect 637 -170 696 -166
rect 534 -250 553 -246
rect -150 -274 -139 -270
rect 46 -270 71 -266
rect -197 -282 -170 -278
rect -197 -323 -187 -282
rect -143 -285 -139 -274
rect -123 -278 -119 -273
rect -27 -277 6 -274
rect -54 -278 6 -277
rect -54 -281 -21 -278
rect -143 -289 -93 -285
rect -123 -307 -119 -289
rect -123 -311 -25 -307
rect -149 -319 -140 -315
rect -29 -319 -25 -311
rect 53 -318 71 -270
rect 146 -266 154 -263
rect 200 -262 204 -258
rect 146 -269 150 -266
rect 154 -315 158 -309
rect 165 -315 169 -309
rect 154 -318 169 -315
rect 505 -266 509 -251
rect 561 -266 565 -250
rect 595 -266 599 -247
rect 637 -258 642 -170
rect 725 -173 729 -163
rect 648 -202 665 -198
rect 651 -207 655 -202
rect 676 -224 681 -193
rect 695 -224 699 -213
rect 703 -214 707 -213
rect 733 -223 737 -213
rect 756 -223 761 -144
rect 791 -156 795 -122
rect 676 -228 726 -224
rect 733 -228 742 -223
rect 747 -228 761 -223
rect 779 -160 795 -156
rect 826 -142 836 -138
rect 779 -188 783 -160
rect 659 -258 663 -247
rect 695 -236 699 -228
rect 733 -236 737 -228
rect 626 -262 652 -258
rect 659 -262 696 -258
rect 492 -270 612 -266
rect -197 -327 -169 -323
rect -197 -352 -187 -327
rect -144 -329 -140 -319
rect -124 -322 -120 -319
rect -83 -325 -47 -321
rect 44 -322 71 -318
rect 173 -321 177 -309
rect 208 -321 212 -282
rect 381 -294 441 -293
rect 626 -294 630 -262
rect 659 -270 663 -262
rect 683 -265 687 -262
rect 725 -265 729 -255
rect 683 -270 729 -265
rect 381 -298 630 -294
rect 651 -295 655 -289
rect -51 -326 -47 -325
rect -144 -333 -103 -329
rect -51 -330 4 -326
rect -149 -348 -136 -344
rect -140 -352 -136 -348
rect -122 -345 -118 -342
rect -82 -348 -71 -344
rect -75 -352 -71 -348
rect -29 -345 -25 -330
rect 53 -344 71 -322
rect 134 -326 218 -321
rect 187 -335 240 -332
rect 187 -338 192 -335
rect 46 -348 71 -344
rect -197 -356 -169 -352
rect -140 -356 -102 -352
rect -75 -356 5 -352
rect -197 -369 -187 -356
rect -82 -365 -69 -361
rect -73 -369 -69 -365
rect -29 -362 -25 -356
rect 53 -361 71 -348
rect 46 -365 71 -361
rect -197 -373 -102 -369
rect -73 -373 6 -369
rect -197 -391 -187 -373
rect -82 -387 -71 -383
rect -197 -395 -102 -391
rect -75 -395 -71 -387
rect -29 -384 -25 -373
rect 53 -383 71 -365
rect 46 -387 71 -383
rect -31 -395 6 -391
rect -197 -413 -187 -395
rect -75 -399 -25 -395
rect -29 -410 -25 -399
rect 53 -406 71 -387
rect 148 -342 207 -338
rect -139 -446 68 -428
rect 148 -430 153 -342
rect 236 -345 240 -335
rect 159 -374 176 -370
rect 162 -379 166 -374
rect 187 -396 192 -365
rect 206 -396 210 -385
rect 214 -386 218 -385
rect 244 -395 248 -385
rect 187 -400 237 -396
rect 244 -400 253 -395
rect 258 -400 284 -395
rect 170 -430 174 -419
rect 206 -408 210 -400
rect 244 -408 248 -400
rect 126 -434 163 -430
rect 170 -434 207 -430
rect -124 -453 -120 -446
rect -72 -453 -68 -446
rect -151 -515 -123 -511
rect -151 -678 -146 -515
rect -116 -527 -112 -493
rect -128 -531 -112 -527
rect -81 -513 -71 -509
rect -128 -559 -124 -531
rect -120 -622 -116 -598
rect -81 -622 -77 -513
rect -64 -520 -60 -493
rect -20 -455 -16 -446
rect 6 -453 10 -446
rect 23 -453 27 -446
rect 45 -453 49 -446
rect -64 -526 -57 -520
rect -12 -524 -8 -495
rect 14 -524 18 -494
rect 31 -524 35 -493
rect 53 -524 57 -493
rect 126 -524 129 -434
rect 170 -442 174 -434
rect 194 -437 198 -434
rect 236 -437 240 -427
rect 194 -442 240 -437
rect 162 -467 166 -461
rect 157 -471 176 -467
rect 162 -504 241 -499
rect -61 -553 -57 -526
rect -31 -528 -19 -524
rect -12 -528 7 -524
rect 14 -528 24 -524
rect 31 -528 46 -524
rect 53 -528 129 -524
rect -53 -618 -49 -592
rect -31 -618 -27 -528
rect -12 -546 -8 -528
rect -17 -550 -8 -546
rect -17 -582 -13 -550
rect 14 -570 18 -528
rect 31 -568 35 -528
rect 53 -530 61 -528
rect 6 -574 18 -570
rect 23 -572 35 -568
rect 57 -570 61 -530
rect 6 -581 10 -574
rect 23 -581 27 -572
rect 45 -574 61 -570
rect 126 -568 129 -528
rect 168 -511 172 -504
rect 187 -511 191 -504
rect 222 -511 226 -504
rect 280 -544 284 -400
rect 381 -543 387 -298
rect 626 -299 630 -298
rect 646 -299 665 -295
rect 756 -307 761 -228
rect 787 -251 791 -227
rect 826 -251 830 -142
rect 843 -149 847 -122
rect 887 -84 891 -75
rect 913 -82 917 -75
rect 930 -82 934 -75
rect 952 -82 956 -75
rect 1064 -82 1068 -75
rect 843 -155 850 -149
rect 895 -153 899 -124
rect 921 -153 925 -123
rect 938 -153 942 -122
rect 960 -153 964 -122
rect 1072 -153 1076 -122
rect 846 -182 850 -155
rect 876 -157 888 -153
rect 895 -157 914 -153
rect 921 -157 931 -153
rect 938 -157 953 -153
rect 960 -157 1065 -153
rect 1072 -157 1093 -153
rect 854 -247 858 -221
rect 876 -247 880 -157
rect 895 -175 899 -157
rect 890 -179 899 -175
rect 890 -211 894 -179
rect 921 -199 925 -157
rect 938 -197 942 -157
rect 960 -159 968 -157
rect 1072 -159 1080 -157
rect 913 -203 925 -199
rect 930 -201 942 -197
rect 964 -199 968 -159
rect 1076 -199 1080 -159
rect 913 -210 917 -203
rect 930 -210 934 -201
rect 952 -203 968 -199
rect 1064 -203 1080 -199
rect 952 -210 956 -203
rect 1064 -210 1068 -203
rect 842 -251 847 -247
rect 854 -251 880 -247
rect 773 -255 780 -251
rect 787 -255 830 -251
rect 787 -269 791 -255
rect 854 -267 858 -251
rect 888 -252 891 -248
rect 779 -273 791 -269
rect 839 -271 858 -267
rect 898 -268 902 -231
rect 911 -250 914 -246
rect 921 -264 925 -230
rect 779 -278 783 -273
rect 839 -278 843 -271
rect 884 -272 902 -268
rect 913 -268 925 -264
rect 884 -277 888 -272
rect 913 -277 917 -268
rect 756 -311 780 -307
rect 787 -315 791 -298
rect 847 -315 851 -298
rect 892 -315 896 -297
rect 921 -315 925 -297
rect 938 -315 942 -230
rect 960 -315 964 -230
rect 1072 -315 1076 -230
rect 778 -325 982 -315
rect 1057 -325 1093 -315
rect 504 -365 688 -359
rect 510 -371 514 -365
rect 530 -371 534 -365
rect 567 -372 571 -365
rect 520 -494 524 -491
rect 553 -376 559 -372
rect 559 -440 563 -432
rect 553 -444 578 -440
rect 663 -383 667 -365
rect 842 -408 1049 -390
rect 1124 -408 1154 -390
rect 752 -419 805 -414
rect 752 -422 757 -419
rect 671 -444 675 -423
rect 713 -426 772 -422
rect 590 -450 660 -444
rect 671 -450 704 -444
rect 671 -459 675 -450
rect 663 -484 667 -479
rect 541 -494 544 -492
rect 520 -497 544 -494
rect 476 -507 511 -503
rect 448 -520 523 -516
rect 413 -534 542 -530
rect 280 -548 381 -544
rect 387 -548 560 -544
rect 280 -549 357 -548
rect 176 -558 180 -551
rect 195 -558 199 -551
rect 230 -558 234 -551
rect 350 -558 355 -555
rect 155 -562 169 -558
rect 181 -562 223 -558
rect 230 -560 355 -558
rect 363 -559 579 -555
rect 230 -561 354 -560
rect 230 -562 353 -561
rect 230 -568 234 -562
rect 586 -563 590 -492
rect 126 -572 188 -568
rect 222 -572 234 -568
rect 541 -567 563 -563
rect 541 -570 545 -567
rect 559 -570 563 -567
rect 578 -567 590 -563
rect 611 -490 690 -484
rect 578 -570 582 -567
rect 45 -581 49 -574
rect 168 -580 176 -577
rect 222 -576 226 -572
rect -65 -622 -60 -618
rect -53 -622 -27 -618
rect -134 -626 -127 -622
rect -120 -626 -77 -622
rect -120 -640 -116 -626
rect -53 -638 -49 -622
rect -19 -623 -16 -619
rect -128 -644 -116 -640
rect -68 -642 -49 -638
rect -9 -639 -5 -602
rect 4 -621 7 -617
rect 14 -635 18 -601
rect -128 -649 -124 -644
rect -68 -649 -64 -642
rect -23 -643 -5 -639
rect 6 -639 18 -635
rect -23 -648 -19 -643
rect 6 -648 10 -639
rect -151 -682 -127 -678
rect -120 -686 -116 -669
rect -60 -686 -56 -669
rect -15 -686 -11 -668
rect 14 -686 18 -668
rect 31 -686 35 -601
rect 53 -686 57 -601
rect 168 -583 172 -580
rect 176 -629 180 -623
rect 187 -629 191 -623
rect 176 -632 191 -629
rect 195 -635 199 -623
rect 230 -635 234 -596
rect 534 -574 541 -570
rect 156 -640 240 -635
rect 510 -638 514 -630
rect 549 -638 553 -600
rect 571 -574 578 -570
rect 586 -638 590 -590
rect 611 -638 615 -490
rect 713 -514 718 -426
rect 801 -429 805 -419
rect 857 -415 861 -408
rect 909 -415 913 -408
rect 724 -458 741 -454
rect 727 -463 731 -458
rect 752 -480 757 -449
rect 771 -480 775 -469
rect 779 -470 783 -469
rect 809 -479 813 -469
rect 830 -477 858 -473
rect 830 -479 835 -477
rect 752 -484 802 -480
rect 809 -484 818 -479
rect 823 -484 835 -479
rect 735 -514 739 -503
rect 771 -492 775 -484
rect 809 -492 813 -484
rect 710 -518 728 -514
rect 735 -518 772 -514
rect 735 -526 739 -518
rect 759 -521 763 -518
rect 801 -521 805 -511
rect 759 -526 805 -521
rect 727 -551 731 -545
rect 722 -555 741 -551
rect 502 -644 615 -638
rect 830 -640 835 -484
rect 865 -489 869 -455
rect 853 -493 869 -489
rect 900 -475 910 -471
rect 853 -521 857 -493
rect 861 -584 865 -560
rect 900 -584 904 -475
rect 917 -482 921 -455
rect 961 -417 965 -408
rect 987 -415 991 -408
rect 1004 -415 1008 -408
rect 1026 -415 1030 -408
rect 1131 -415 1135 -408
rect 917 -488 924 -482
rect 969 -486 973 -457
rect 995 -486 999 -456
rect 1012 -486 1016 -455
rect 1034 -486 1038 -455
rect 1139 -486 1143 -455
rect 920 -515 924 -488
rect 950 -490 962 -486
rect 969 -490 988 -486
rect 995 -490 1005 -486
rect 1012 -490 1027 -486
rect 1034 -490 1132 -486
rect 1139 -490 1160 -486
rect 928 -580 932 -554
rect 950 -580 954 -490
rect 969 -508 973 -490
rect 964 -512 973 -508
rect 964 -544 968 -512
rect 995 -532 999 -490
rect 1012 -530 1016 -490
rect 1034 -492 1042 -490
rect 1139 -492 1147 -490
rect 987 -536 999 -532
rect 1004 -534 1016 -530
rect 1038 -532 1042 -492
rect 1143 -532 1147 -492
rect 987 -543 991 -536
rect 1004 -543 1008 -534
rect 1026 -536 1042 -532
rect 1131 -536 1147 -532
rect 1026 -543 1030 -536
rect 1131 -543 1135 -536
rect 916 -584 921 -580
rect 928 -584 954 -580
rect 847 -588 854 -584
rect 861 -588 904 -584
rect 861 -602 865 -588
rect 928 -600 932 -584
rect 962 -585 965 -581
rect 853 -606 865 -602
rect 913 -604 932 -600
rect 972 -601 976 -564
rect 985 -583 988 -579
rect 995 -597 999 -563
rect 853 -611 857 -606
rect 913 -611 917 -604
rect 958 -605 976 -601
rect 987 -601 999 -597
rect 958 -610 962 -605
rect 987 -610 991 -601
rect 830 -644 854 -640
rect 861 -648 865 -631
rect 921 -648 925 -631
rect 966 -648 970 -630
rect 995 -648 999 -630
rect 1012 -648 1016 -563
rect 1034 -648 1038 -563
rect 1139 -648 1143 -563
rect 852 -658 1056 -648
rect 1124 -658 1160 -648
rect 500 -671 696 -665
rect 509 -678 513 -671
rect 535 -678 539 -671
rect 571 -678 575 -671
rect 609 -677 613 -671
rect -129 -696 75 -686
rect -119 -725 88 -707
rect -104 -732 -100 -725
rect -52 -732 -48 -725
rect -131 -794 -103 -790
rect -131 -857 -126 -794
rect -96 -806 -92 -772
rect -137 -861 -126 -857
rect -131 -885 -126 -861
rect -108 -810 -92 -806
rect -61 -792 -51 -788
rect -108 -838 -104 -810
rect -132 -890 -126 -885
rect -131 -957 -126 -890
rect -100 -901 -96 -877
rect -61 -901 -57 -792
rect -44 -799 -40 -772
rect 0 -734 4 -725
rect 26 -732 30 -725
rect 43 -732 47 -725
rect 65 -732 69 -725
rect 187 -764 240 -759
rect 187 -767 192 -764
rect -44 -805 -37 -799
rect 8 -803 12 -774
rect 34 -803 38 -773
rect 51 -803 55 -772
rect 73 -803 77 -772
rect 148 -771 207 -767
rect -41 -832 -37 -805
rect -11 -807 1 -803
rect 8 -807 27 -803
rect 34 -807 44 -803
rect 51 -807 66 -803
rect 73 -807 107 -803
rect -33 -897 -29 -871
rect -11 -897 -7 -807
rect 8 -825 12 -807
rect 3 -829 12 -825
rect 3 -861 7 -829
rect 34 -849 38 -807
rect 51 -847 55 -807
rect 73 -809 81 -807
rect 26 -853 38 -849
rect 43 -851 55 -847
rect 77 -849 81 -809
rect 26 -860 30 -853
rect 43 -860 47 -851
rect 65 -853 81 -849
rect 65 -860 69 -853
rect 148 -859 153 -771
rect 236 -774 240 -764
rect 159 -803 176 -799
rect 162 -808 166 -803
rect 187 -825 192 -794
rect 206 -825 210 -814
rect 214 -815 218 -814
rect 244 -824 248 -814
rect 265 -824 269 -823
rect 187 -829 237 -825
rect 244 -829 253 -824
rect 258 -829 269 -824
rect 170 -859 174 -848
rect 206 -837 210 -829
rect 244 -837 248 -829
rect -45 -901 -40 -897
rect -33 -901 -7 -897
rect -114 -905 -107 -901
rect -100 -905 -57 -901
rect -100 -919 -96 -905
rect -33 -917 -29 -901
rect 1 -902 4 -898
rect -108 -923 -96 -919
rect -48 -921 -29 -917
rect 11 -918 15 -881
rect 24 -900 27 -896
rect 34 -914 38 -880
rect -108 -928 -104 -923
rect -48 -928 -44 -921
rect -3 -922 15 -918
rect 26 -918 38 -914
rect -3 -927 1 -922
rect 26 -927 30 -918
rect -131 -961 -107 -957
rect -100 -965 -96 -948
rect -40 -965 -36 -948
rect 5 -965 9 -947
rect 34 -965 38 -947
rect 51 -965 55 -880
rect 73 -965 77 -880
rect 126 -863 163 -859
rect 170 -863 207 -859
rect -109 -975 95 -965
rect 126 -997 129 -863
rect 170 -871 174 -863
rect 194 -866 198 -863
rect 236 -866 240 -856
rect 194 -871 240 -866
rect 162 -896 166 -890
rect 157 -900 176 -896
rect 162 -933 241 -928
rect 168 -940 172 -933
rect 187 -940 191 -933
rect 222 -940 226 -933
rect 264 -955 269 -829
rect 521 -683 527 -678
rect 557 -682 563 -678
rect 563 -764 567 -758
rect 563 -768 582 -764
rect 594 -682 601 -677
rect 601 -742 605 -731
rect 601 -746 619 -742
rect 527 -848 531 -838
rect 545 -848 549 -838
rect 475 -855 509 -848
rect 526 -852 549 -848
rect 590 -849 594 -837
rect 619 -849 623 -836
rect 590 -853 623 -849
rect 652 -677 656 -671
rect 448 -874 527 -867
rect 413 -892 545 -885
rect 387 -913 563 -906
rect 363 -935 582 -928
rect 264 -962 326 -955
rect 333 -962 601 -955
rect 627 -962 631 -836
rect 660 -962 664 -717
rect 835 -836 1042 -818
rect 1124 -836 1154 -818
rect 850 -843 854 -836
rect 902 -843 906 -836
rect 823 -905 851 -901
rect 743 -936 796 -931
rect 743 -939 748 -936
rect 704 -943 763 -939
rect 176 -987 180 -980
rect 195 -987 199 -980
rect 230 -987 234 -980
rect 627 -966 653 -962
rect 660 -966 695 -962
rect 291 -987 294 -984
rect 155 -991 169 -987
rect 181 -991 223 -987
rect 230 -991 294 -987
rect 299 -991 619 -984
rect 230 -997 234 -991
rect 20 -1001 188 -997
rect 222 -1001 234 -997
rect 20 -1002 150 -1001
rect -121 -1078 -103 -1059
rect 20 -1066 25 -1002
rect 168 -1009 176 -1006
rect 222 -1005 226 -1001
rect 168 -1012 172 -1009
rect -25 -1070 25 -1066
rect 137 -1070 147 -1052
rect 176 -1058 180 -1052
rect 187 -1058 191 -1052
rect 176 -1061 191 -1058
rect 627 -1008 631 -966
rect 195 -1064 199 -1052
rect 230 -1064 234 -1025
rect 156 -1069 240 -1064
rect -56 -1074 -19 -1070
rect -121 -1082 -96 -1078
rect -121 -1100 -103 -1082
rect -25 -1092 -21 -1081
rect 21 -1078 25 -1070
rect 52 -1074 147 -1070
rect 21 -1082 32 -1078
rect 137 -1092 147 -1074
rect -56 -1096 23 -1092
rect 52 -1096 147 -1092
rect -121 -1104 -96 -1100
rect -121 -1117 -103 -1104
rect -25 -1109 -21 -1103
rect 19 -1100 23 -1096
rect 19 -1104 32 -1100
rect 137 -1109 147 -1096
rect 521 -1088 527 -1083
rect 509 -1106 513 -1088
rect 539 -1013 563 -1009
rect 539 -1088 545 -1084
rect 539 -1089 549 -1088
rect 553 -1106 557 -1088
rect 575 -1013 601 -1009
rect 575 -1088 582 -1084
rect 613 -1012 633 -1008
rect 660 -1068 664 -966
rect 704 -1031 709 -943
rect 792 -946 796 -936
rect 715 -975 732 -971
rect 718 -980 722 -975
rect 743 -997 748 -966
rect 762 -997 766 -986
rect 770 -987 774 -986
rect 800 -996 804 -986
rect 823 -996 828 -905
rect 858 -917 862 -883
rect 846 -921 862 -917
rect 893 -903 903 -899
rect 846 -949 850 -921
rect 743 -1001 793 -997
rect 800 -1001 809 -996
rect 814 -1001 828 -996
rect 726 -1031 730 -1020
rect 762 -1009 766 -1001
rect 800 -1009 804 -1001
rect 613 -1088 619 -1084
rect 590 -1106 594 -1088
rect 627 -1106 631 -1088
rect 696 -1035 719 -1031
rect 726 -1035 763 -1031
rect 652 -1106 656 -1088
rect -55 -1113 25 -1109
rect 52 -1113 90 -1109
rect 119 -1113 147 -1109
rect 486 -1112 669 -1106
rect -121 -1121 -96 -1117
rect -121 -1143 -103 -1121
rect -25 -1135 -21 -1120
rect 21 -1117 25 -1113
rect 21 -1121 32 -1117
rect 68 -1123 72 -1120
rect 86 -1117 90 -1113
rect 86 -1121 99 -1117
rect -54 -1139 1 -1135
rect 53 -1136 94 -1132
rect -3 -1140 1 -1139
rect -121 -1147 -94 -1143
rect -3 -1144 33 -1140
rect 70 -1146 74 -1143
rect 90 -1146 94 -1136
rect 137 -1138 147 -1113
rect 696 -1127 701 -1035
rect 726 -1043 730 -1035
rect 750 -1038 754 -1035
rect 792 -1038 796 -1028
rect 750 -1043 796 -1038
rect 718 -1068 722 -1062
rect 823 -1068 828 -1001
rect 854 -1012 858 -988
rect 893 -1012 897 -903
rect 910 -910 914 -883
rect 954 -845 958 -836
rect 980 -843 984 -836
rect 997 -843 1001 -836
rect 1019 -843 1023 -836
rect 1131 -843 1135 -836
rect 910 -916 917 -910
rect 962 -914 966 -885
rect 988 -914 992 -884
rect 1005 -914 1009 -883
rect 1027 -914 1031 -883
rect 1139 -914 1143 -883
rect 913 -943 917 -916
rect 943 -918 955 -914
rect 962 -918 981 -914
rect 988 -918 998 -914
rect 1005 -918 1020 -914
rect 1027 -918 1132 -914
rect 1139 -918 1160 -914
rect 921 -1008 925 -982
rect 943 -1008 947 -918
rect 962 -936 966 -918
rect 957 -940 966 -936
rect 957 -972 961 -940
rect 988 -960 992 -918
rect 1005 -958 1009 -918
rect 1027 -920 1035 -918
rect 1139 -920 1147 -918
rect 980 -964 992 -960
rect 997 -962 1009 -958
rect 1031 -960 1035 -920
rect 1143 -960 1147 -920
rect 980 -971 984 -964
rect 997 -971 1001 -962
rect 1019 -964 1035 -960
rect 1131 -964 1147 -960
rect 1019 -971 1023 -964
rect 1131 -971 1135 -964
rect 909 -1012 914 -1008
rect 921 -1012 947 -1008
rect 840 -1016 847 -1012
rect 854 -1016 897 -1012
rect 854 -1030 858 -1016
rect 921 -1028 925 -1012
rect 955 -1013 958 -1009
rect 846 -1034 858 -1030
rect 906 -1032 925 -1028
rect 965 -1029 969 -992
rect 978 -1011 981 -1007
rect 988 -1025 992 -991
rect 846 -1039 850 -1034
rect 906 -1039 910 -1032
rect 951 -1033 969 -1029
rect 980 -1029 992 -1025
rect 951 -1038 955 -1033
rect 980 -1038 984 -1029
rect 713 -1072 732 -1068
rect 823 -1072 847 -1068
rect 854 -1076 858 -1059
rect 914 -1076 918 -1059
rect 959 -1076 963 -1058
rect 988 -1076 992 -1058
rect 1005 -1076 1009 -991
rect 1027 -1076 1031 -991
rect 1139 -1076 1143 -991
rect 845 -1086 1049 -1076
rect 1124 -1086 1160 -1076
rect 119 -1142 147 -1138
rect -121 -1195 -103 -1147
rect -25 -1154 -21 -1146
rect 90 -1150 99 -1146
rect -25 -1158 73 -1154
rect 69 -1176 73 -1158
rect 43 -1180 93 -1176
rect -29 -1187 4 -1184
rect -56 -1188 4 -1187
rect -56 -1191 -23 -1188
rect 69 -1192 73 -1187
rect 89 -1191 93 -1180
rect 137 -1183 147 -1142
rect 493 -1146 700 -1142
rect 120 -1187 147 -1183
rect -121 -1199 -96 -1195
rect 89 -1195 100 -1191
rect -121 -1247 -103 -1199
rect -40 -1204 -36 -1198
rect -40 -1208 77 -1204
rect -56 -1243 -18 -1239
rect 73 -1243 77 -1208
rect 137 -1243 147 -1187
rect -121 -1251 -96 -1247
rect -121 -1266 -103 -1251
rect -38 -1273 -34 -1250
rect -22 -1251 -18 -1243
rect 49 -1247 95 -1243
rect 120 -1247 147 -1243
rect -22 -1255 10 -1251
rect 73 -1261 77 -1254
rect 91 -1251 95 -1247
rect 91 -1255 100 -1251
rect 129 -1273 133 -1254
rect 137 -1256 147 -1247
rect 499 -1155 503 -1146
rect 526 -1155 530 -1146
rect 562 -1155 566 -1146
rect 597 -1155 601 -1146
rect 634 -1155 638 -1146
rect -38 -1278 133 -1273
rect 29 -1280 33 -1278
rect 57 -1279 62 -1278
rect 190 -1293 243 -1288
rect 190 -1296 195 -1293
rect 151 -1300 210 -1296
rect -121 -1335 86 -1317
rect -106 -1342 -102 -1335
rect -54 -1342 -50 -1335
rect -133 -1404 -105 -1400
rect -133 -1467 -128 -1404
rect -98 -1416 -94 -1382
rect -135 -1471 -128 -1467
rect -133 -1495 -128 -1471
rect -110 -1420 -94 -1416
rect -63 -1402 -53 -1398
rect -110 -1448 -106 -1420
rect -134 -1500 -128 -1495
rect -133 -1567 -128 -1500
rect -102 -1511 -98 -1487
rect -63 -1511 -59 -1402
rect -46 -1409 -42 -1382
rect -2 -1344 2 -1335
rect 24 -1342 28 -1335
rect 41 -1342 45 -1335
rect 63 -1342 67 -1335
rect -46 -1415 -39 -1409
rect 6 -1413 10 -1384
rect 32 -1413 36 -1383
rect 49 -1413 53 -1382
rect 71 -1413 75 -1382
rect 151 -1388 156 -1300
rect 239 -1303 243 -1293
rect 162 -1332 179 -1328
rect 165 -1337 169 -1332
rect 190 -1354 195 -1323
rect 209 -1354 213 -1343
rect 217 -1344 221 -1343
rect 247 -1353 251 -1343
rect 190 -1358 240 -1354
rect 247 -1358 256 -1353
rect 261 -1358 270 -1353
rect 511 -1159 518 -1155
rect 511 -1354 518 -1351
rect 173 -1388 177 -1377
rect 209 -1366 213 -1358
rect 247 -1366 251 -1358
rect 129 -1392 166 -1388
rect 173 -1392 210 -1388
rect -43 -1442 -39 -1415
rect -13 -1417 -1 -1413
rect 6 -1417 25 -1413
rect 32 -1417 42 -1413
rect 49 -1417 64 -1413
rect 71 -1417 109 -1413
rect -35 -1507 -31 -1481
rect -13 -1507 -9 -1417
rect 6 -1435 10 -1417
rect 1 -1439 10 -1435
rect 1 -1471 5 -1439
rect 32 -1459 36 -1417
rect 49 -1457 53 -1417
rect 71 -1419 79 -1417
rect 24 -1463 36 -1459
rect 41 -1461 53 -1457
rect 75 -1459 79 -1419
rect 24 -1470 28 -1463
rect 41 -1470 45 -1461
rect 63 -1463 79 -1459
rect 63 -1470 67 -1463
rect -47 -1511 -42 -1507
rect -35 -1511 -9 -1507
rect -116 -1515 -109 -1511
rect -102 -1515 -59 -1511
rect -102 -1529 -98 -1515
rect -35 -1527 -31 -1511
rect -1 -1512 2 -1508
rect -110 -1533 -98 -1529
rect -50 -1531 -31 -1527
rect 9 -1528 13 -1491
rect 22 -1510 25 -1506
rect 32 -1524 36 -1490
rect -110 -1538 -106 -1533
rect -50 -1538 -46 -1531
rect -5 -1532 13 -1528
rect 24 -1528 36 -1524
rect -5 -1537 -1 -1532
rect 24 -1537 28 -1528
rect -133 -1571 -109 -1567
rect -102 -1575 -98 -1558
rect -42 -1575 -38 -1558
rect 3 -1575 7 -1557
rect 32 -1575 36 -1557
rect 49 -1575 53 -1490
rect 71 -1575 75 -1490
rect 129 -1526 132 -1392
rect 173 -1400 177 -1392
rect 197 -1395 201 -1392
rect 239 -1395 243 -1385
rect 197 -1400 243 -1395
rect 165 -1425 169 -1419
rect 160 -1429 179 -1425
rect 165 -1462 244 -1457
rect 171 -1469 175 -1462
rect 190 -1469 194 -1462
rect 225 -1469 229 -1462
rect 271 -1498 275 -1358
rect 518 -1358 522 -1355
rect 536 -1358 540 -1355
rect 518 -1362 540 -1358
rect 548 -1159 554 -1155
rect 544 -1357 548 -1355
rect 583 -1159 589 -1155
rect 583 -1355 607 -1351
rect 619 -1160 626 -1155
rect 619 -1355 645 -1351
rect 681 -1169 685 -1146
rect 571 -1357 575 -1355
rect 544 -1362 575 -1357
rect 475 -1399 499 -1394
rect 653 -1402 657 -1355
rect 689 -1400 693 -1209
rect 728 -1268 935 -1250
rect 1017 -1268 1047 -1250
rect 743 -1275 747 -1268
rect 795 -1275 799 -1268
rect 716 -1337 744 -1333
rect 716 -1400 721 -1337
rect 751 -1349 755 -1315
rect 653 -1403 680 -1402
rect 447 -1413 518 -1408
rect 653 -1409 681 -1403
rect 689 -1404 721 -1400
rect 412 -1430 536 -1425
rect 386 -1444 554 -1439
rect 362 -1460 571 -1455
rect 332 -1473 589 -1468
rect 299 -1490 607 -1485
rect 271 -1499 474 -1498
rect 271 -1504 626 -1499
rect 271 -1505 504 -1504
rect 179 -1516 183 -1509
rect 198 -1516 202 -1509
rect 233 -1516 237 -1509
rect 455 -1516 645 -1515
rect 158 -1520 172 -1516
rect 184 -1520 226 -1516
rect 233 -1520 645 -1516
rect 233 -1526 237 -1520
rect 129 -1530 191 -1526
rect 225 -1530 237 -1526
rect -111 -1585 93 -1575
rect 47 -1618 65 -1599
rect 143 -1606 147 -1530
rect 171 -1538 179 -1535
rect 225 -1534 229 -1530
rect 171 -1541 175 -1538
rect 179 -1587 183 -1581
rect 190 -1587 194 -1581
rect 179 -1590 194 -1587
rect 198 -1593 202 -1581
rect 233 -1593 237 -1554
rect 159 -1598 243 -1593
rect 143 -1610 193 -1606
rect 305 -1610 315 -1592
rect 112 -1614 149 -1610
rect 47 -1622 72 -1618
rect 47 -1640 65 -1622
rect 143 -1632 147 -1621
rect 189 -1618 193 -1610
rect 220 -1614 315 -1610
rect 189 -1622 200 -1618
rect 305 -1632 315 -1614
rect 112 -1636 191 -1632
rect 220 -1636 315 -1632
rect 47 -1644 72 -1640
rect 47 -1657 65 -1644
rect 143 -1649 147 -1643
rect 187 -1640 191 -1636
rect 187 -1644 200 -1640
rect 305 -1649 315 -1636
rect 499 -1637 503 -1632
rect 511 -1632 518 -1630
rect 530 -1537 554 -1532
rect 530 -1632 536 -1628
rect 566 -1536 589 -1532
rect 566 -1632 571 -1628
rect 601 -1536 626 -1532
rect 601 -1632 607 -1628
rect 653 -1598 657 -1409
rect 645 -1601 657 -1598
rect 645 -1612 649 -1601
rect 689 -1612 693 -1404
rect 716 -1428 721 -1404
rect 739 -1353 755 -1349
rect 786 -1335 796 -1331
rect 739 -1381 743 -1353
rect 715 -1433 721 -1428
rect 716 -1500 721 -1433
rect 747 -1444 751 -1420
rect 786 -1444 790 -1335
rect 803 -1342 807 -1315
rect 847 -1277 851 -1268
rect 873 -1275 877 -1268
rect 890 -1275 894 -1268
rect 912 -1275 916 -1268
rect 1024 -1275 1028 -1268
rect 803 -1348 810 -1342
rect 855 -1346 859 -1317
rect 881 -1346 885 -1316
rect 898 -1346 902 -1315
rect 920 -1346 924 -1315
rect 1032 -1346 1036 -1315
rect 806 -1375 810 -1348
rect 836 -1350 848 -1346
rect 855 -1350 874 -1346
rect 881 -1350 891 -1346
rect 898 -1350 913 -1346
rect 920 -1350 1025 -1346
rect 1032 -1350 1053 -1346
rect 814 -1440 818 -1414
rect 836 -1440 840 -1350
rect 855 -1368 859 -1350
rect 850 -1372 859 -1368
rect 850 -1404 854 -1372
rect 881 -1392 885 -1350
rect 898 -1390 902 -1350
rect 920 -1352 928 -1350
rect 1032 -1352 1040 -1350
rect 873 -1396 885 -1392
rect 890 -1394 902 -1390
rect 924 -1392 928 -1352
rect 1036 -1392 1040 -1352
rect 873 -1403 877 -1396
rect 890 -1403 894 -1394
rect 912 -1396 928 -1392
rect 1024 -1396 1040 -1392
rect 912 -1403 916 -1396
rect 1024 -1403 1028 -1396
rect 802 -1444 807 -1440
rect 814 -1444 840 -1440
rect 733 -1448 740 -1444
rect 747 -1448 790 -1444
rect 747 -1462 751 -1448
rect 814 -1460 818 -1444
rect 848 -1445 851 -1441
rect 739 -1466 751 -1462
rect 799 -1464 818 -1460
rect 858 -1461 862 -1424
rect 871 -1443 874 -1439
rect 881 -1457 885 -1423
rect 739 -1471 743 -1466
rect 799 -1471 803 -1464
rect 844 -1465 862 -1461
rect 873 -1461 885 -1457
rect 844 -1470 848 -1465
rect 873 -1470 877 -1461
rect 716 -1504 740 -1500
rect 747 -1508 751 -1491
rect 807 -1508 811 -1491
rect 852 -1508 856 -1490
rect 881 -1508 885 -1490
rect 898 -1508 902 -1423
rect 920 -1508 924 -1423
rect 1032 -1508 1036 -1423
rect 738 -1518 942 -1508
rect 1017 -1518 1053 -1508
rect 638 -1632 645 -1628
rect 507 -1634 522 -1632
rect 544 -1637 548 -1632
rect 579 -1637 583 -1632
rect 615 -1637 619 -1632
rect 653 -1637 657 -1632
rect 681 -1637 685 -1632
rect 488 -1641 694 -1637
rect 113 -1653 193 -1649
rect 220 -1653 258 -1649
rect 287 -1653 315 -1649
rect 47 -1661 72 -1657
rect 47 -1683 65 -1661
rect 143 -1675 147 -1660
rect 189 -1657 193 -1653
rect 189 -1661 200 -1657
rect 236 -1663 240 -1660
rect 254 -1657 258 -1653
rect 254 -1661 267 -1657
rect 114 -1679 169 -1675
rect 221 -1676 262 -1672
rect 165 -1680 169 -1679
rect 47 -1687 74 -1683
rect 165 -1684 201 -1680
rect 238 -1686 242 -1683
rect 258 -1686 262 -1676
rect 305 -1678 315 -1653
rect 287 -1682 315 -1678
rect 47 -1735 65 -1687
rect 143 -1694 147 -1686
rect 258 -1690 267 -1686
rect 143 -1698 241 -1694
rect 237 -1716 241 -1698
rect 211 -1720 261 -1716
rect 139 -1727 172 -1724
rect 112 -1728 172 -1727
rect 112 -1731 145 -1728
rect 237 -1732 241 -1727
rect 257 -1731 261 -1720
rect 305 -1723 315 -1682
rect 288 -1727 315 -1723
rect 47 -1739 72 -1735
rect 257 -1735 268 -1731
rect 47 -1787 65 -1739
rect 128 -1744 132 -1738
rect 128 -1748 245 -1744
rect 112 -1783 150 -1779
rect 241 -1783 245 -1748
rect 305 -1783 315 -1727
rect 47 -1791 72 -1787
rect 47 -1806 65 -1791
rect 130 -1813 134 -1790
rect 146 -1791 150 -1783
rect 217 -1787 263 -1783
rect 288 -1787 315 -1783
rect 146 -1795 178 -1791
rect 241 -1801 245 -1794
rect 259 -1791 263 -1787
rect 259 -1795 268 -1791
rect 297 -1813 301 -1794
rect 305 -1796 315 -1787
rect 130 -1818 301 -1813
rect 197 -1820 201 -1818
rect 225 -1819 230 -1818
<< metal2 >>
rect 375 111 379 115
rect 74 90 78 94
rect 377 88 381 92
rect 76 67 80 71
rect 728 57 762 61
rect 474 19 691 24
rect 728 -2 733 57
rect 758 53 762 57
rect 723 -7 733 -2
rect 202 -13 236 -9
rect 83 -46 89 -43
rect 89 -51 165 -46
rect -98 -100 -94 -96
rect -75 -98 -71 -94
rect 85 -244 89 -51
rect 202 -72 207 -13
rect 232 -17 236 -13
rect 197 -77 207 -72
rect 192 -89 197 -77
rect 231 -81 236 -17
rect 404 -14 620 -8
rect 404 -80 411 -14
rect 718 -19 723 -7
rect 757 -11 762 53
rect 901 44 905 48
rect 924 46 928 50
rect 713 -155 747 -151
rect 634 -193 676 -188
rect 713 -214 718 -155
rect 743 -159 747 -155
rect 708 -219 718 -214
rect 703 -231 708 -219
rect 742 -223 747 -159
rect 85 -249 128 -244
rect 154 -261 159 -249
rect 891 -252 895 -248
rect 914 -250 918 -246
rect -124 -326 -120 -322
rect -122 -349 -118 -345
rect 107 -365 187 -360
rect 107 -411 111 -365
rect 224 -369 229 -332
rect 253 -369 258 -332
rect 224 -373 258 -369
rect 224 -386 229 -373
rect 219 -391 229 -386
rect 214 -403 219 -391
rect 253 -395 258 -373
rect -24 -416 111 -411
rect 107 -558 111 -416
rect 789 -411 823 -407
rect 709 -449 752 -444
rect 789 -470 794 -411
rect 819 -415 823 -411
rect 784 -475 794 -470
rect 779 -487 784 -475
rect 818 -479 823 -415
rect 107 -563 150 -558
rect 176 -575 181 -563
rect -16 -623 -12 -619
rect 7 -621 11 -617
rect 705 -653 709 -518
rect 965 -585 969 -581
rect 988 -583 992 -579
rect 326 -658 709 -653
rect 224 -756 258 -752
rect 107 -794 187 -789
rect 107 -802 111 -794
rect 4 -902 8 -898
rect 27 -900 31 -896
rect 107 -987 111 -807
rect 224 -815 229 -756
rect 254 -760 258 -756
rect 219 -820 229 -815
rect 214 -832 219 -820
rect 253 -824 258 -760
rect 326 -955 333 -658
rect 780 -928 814 -924
rect 700 -966 743 -961
rect 107 -992 150 -987
rect 780 -987 785 -928
rect 810 -932 814 -928
rect 176 -1004 181 -992
rect 775 -992 785 -987
rect 770 -1004 775 -992
rect 809 -996 814 -932
rect 958 -1013 962 -1009
rect 981 -1011 985 -1007
rect 68 -1120 72 -1116
rect 270 -1132 696 -1127
rect 270 -1134 276 -1132
rect 70 -1143 74 -1139
rect 227 -1285 261 -1281
rect 110 -1318 115 -1317
rect 110 -1323 190 -1318
rect 110 -1412 114 -1323
rect 227 -1344 232 -1285
rect 257 -1289 261 -1285
rect 222 -1349 232 -1344
rect 217 -1361 222 -1349
rect 256 -1353 261 -1289
rect 270 -1353 275 -1134
rect 2 -1512 6 -1508
rect 25 -1510 29 -1506
rect 110 -1516 114 -1418
rect 851 -1445 855 -1441
rect 874 -1443 878 -1439
rect 110 -1521 153 -1516
rect 179 -1533 184 -1521
rect 236 -1660 240 -1656
rect 238 -1683 242 -1679
<< m123contact >>
rect 468 19 474 24
rect 691 19 696 24
rect 718 -7 723 -2
rect 83 -51 89 -46
rect 165 -51 170 -46
rect 192 -77 197 -72
rect 620 -15 625 -7
rect 757 -16 762 -11
rect 718 -24 723 -19
rect 231 -86 236 -81
rect 403 -86 411 -80
rect 192 -94 197 -89
rect 470 -137 475 -132
rect 441 -176 448 -170
rect 628 -193 634 -187
rect 676 -193 681 -188
rect 703 -219 708 -214
rect 742 -228 747 -223
rect 703 -236 708 -231
rect 128 -249 133 -244
rect 154 -249 159 -244
rect 406 -249 412 -243
rect 154 -266 159 -261
rect 187 -365 192 -360
rect -30 -417 -24 -410
rect 214 -391 219 -386
rect 253 -400 258 -395
rect 214 -408 219 -403
rect 704 -450 709 -444
rect 752 -449 757 -444
rect 779 -475 784 -470
rect 818 -484 823 -479
rect 779 -492 784 -487
rect 469 -508 476 -502
rect 441 -521 448 -515
rect 705 -518 710 -513
rect 406 -535 413 -529
rect 381 -548 387 -543
rect 150 -563 155 -558
rect 176 -563 181 -558
rect 355 -560 363 -555
rect 176 -580 181 -575
rect 187 -794 192 -789
rect 107 -807 112 -802
rect 214 -820 219 -815
rect 253 -829 258 -824
rect 214 -837 219 -832
rect 469 -855 475 -848
rect 442 -874 448 -867
rect 407 -892 413 -885
rect 381 -913 387 -906
rect 356 -935 363 -928
rect 326 -962 333 -955
rect 695 -966 700 -961
rect 743 -966 748 -961
rect 150 -992 155 -987
rect 176 -992 181 -987
rect 294 -991 299 -984
rect 176 -1009 181 -1004
rect 770 -992 775 -987
rect 809 -1001 814 -996
rect 770 -1009 775 -1004
rect 696 -1132 701 -1127
rect 190 -1323 195 -1318
rect 217 -1349 222 -1344
rect 256 -1358 261 -1353
rect 270 -1358 275 -1353
rect 217 -1366 222 -1361
rect 470 -1399 475 -1394
rect 109 -1418 115 -1412
rect 442 -1413 447 -1408
rect 407 -1430 412 -1425
rect 381 -1444 386 -1439
rect 356 -1460 362 -1455
rect 326 -1473 332 -1468
rect 294 -1490 299 -1485
rect 153 -1521 158 -1516
rect 179 -1521 184 -1516
rect 179 -1538 184 -1533
<< metal3 >>
rect 470 -132 474 19
rect 407 -529 412 -249
rect 442 -515 447 -176
rect 470 -502 475 -137
rect 356 -928 363 -560
rect 381 -906 387 -548
rect 407 -885 412 -535
rect 442 -867 447 -521
rect 470 -644 475 -508
rect 470 -667 476 -644
rect 470 -848 475 -667
rect 294 -1099 299 -991
rect 294 -1141 300 -1099
rect 294 -1485 299 -1141
rect 326 -1468 332 -962
rect 356 -1104 362 -935
rect 355 -1117 362 -1104
rect 381 -1100 386 -913
rect 407 -1099 412 -892
rect 355 -1140 361 -1117
rect 355 -1146 362 -1140
rect 356 -1455 362 -1146
rect 381 -1142 387 -1100
rect 406 -1141 412 -1099
rect 381 -1439 386 -1142
rect 407 -1425 412 -1141
rect 442 -1100 447 -874
rect 442 -1142 448 -1100
rect 470 -1101 475 -855
rect 442 -1408 447 -1142
rect 470 -1143 476 -1101
rect 470 -1394 475 -1143
<< labels >>
rlabel metal1 138 -432 141 -431 1 b2
rlabel metal2 118 -364 121 -363 1 a2
rlabel metal1 160 -470 165 -469 1 gnd2
rlabel metal1 163 -372 168 -371 1 vdd2
rlabel metal1 110 -119 115 -117 1 b1
rlabel metal2 104 -50 109 -48 1 a1
rlabel metal1 141 -59 147 -57 1 vdd11
rlabel metal1 138 -156 144 -154 1 gnd11
rlabel metal1 254 -84 258 -83 1 p1
rlabel metal1 266 -397 276 -396 1 p2
rlabel metal1 246 -246 246 -246 1 g1
rlabel metal1 186 -325 192 -323 1 gnd1
rlabel metal1 176 -188 182 -186 5 vdd1
rlabel metal1 270 -561 280 -560 1 g2
rlabel metal1 178 -501 183 -500 1 vdd22
rlabel metal1 182 -637 187 -636 1 gnd22
rlabel metal1 614 -134 618 -132 1 c1
rlabel metal1 538 -269 538 -269 1 gndc1
rlabel metal1 527 -31 532 -29 1 vddc1
rlabel metal1 666 10 666 10 1 vdds1
rlabel metal1 764 -14 765 -14 1 s1
rlabel metal1 669 -83 669 -83 1 gnds1
rlabel metal1 654 -201 654 -201 1 vdds2
rlabel metal1 653 -297 653 -297 1 gnds2
rlabel metal1 553 -361 557 -360 1 vddc2
rlabel metal1 517 -642 520 -641 1 gndc2
rlabel metal1 477 -960 483 -957 1 p3
rlabel metal1 682 -964 690 -962 1 c3
rlabel metal1 478 -989 484 -986 1 g3
rlabel metal1 543 -668 551 -667 1 vddc3
rlabel metal1 580 -1110 582 -1109 1 gndc3
rlabel metal1 182 -1066 187 -1065 1 gnd33
rlabel metal1 178 -930 183 -929 1 vdd33
rlabel metal2 118 -793 121 -792 1 a3
rlabel metal1 138 -861 141 -860 1 b3
rlabel metal1 160 -899 165 -898 1 gnd3
rlabel metal1 163 -801 168 -800 1 vdd3
rlabel metal1 735 -553 735 -553 1 gnds3
rlabel metal1 732 -457 732 -457 1 vdds3
rlabel metal1 700 -447 703 -446 1 c2
rlabel metal1 827 -481 827 -481 1 s3
rlabel metal1 566 -1640 566 -1640 1 gndc4
rlabel metal1 622 -1143 622 -1143 1 vddc4
rlabel metal1 700 -1402 700 -1402 1 c4
rlabel metal1 476 -1519 477 -1518 1 g4
rlabel metal1 475 -1503 476 -1502 1 p4
rlabel metal1 196 -1595 198 -1594 1 gnd44
rlabel metal1 168 -1330 170 -1329 1 vdd4
rlabel metal1 182 -1460 184 -1459 1 vdd44
rlabel metal1 165 -1428 167 -1427 1 gnd4
rlabel metal1 134 -1391 137 -1390 1 b4
rlabel metal1 819 -998 819 -998 1 s4
rlabel metal1 720 -973 720 -973 1 vdds4
rlabel metal1 717 -1070 717 -1070 1 gnds4
rlabel metal1 750 -225 750 -225 1 s2
rlabel metal1 785 43 785 43 1 clk
rlabel metal1 854 47 854 47 1 clk
rlabel metal1 900 46 900 46 1 clk
rlabel metal1 922 47 922 47 1 clk
rlabel metal1 988 141 988 141 1 s1o
rlabel metal1 867 231 867 231 1 vdd
rlabel metal1 959 -25 959 -25 1 gnd
rlabel metal1 949 -321 949 -321 1 gnd
rlabel metal1 857 -65 857 -65 1 vdd
rlabel metal1 912 -249 912 -249 1 clk
rlabel metal1 890 -250 890 -250 1 clk
rlabel metal1 844 -249 844 -249 1 clk
rlabel metal1 775 -253 775 -253 1 clk
rlabel metal1 978 -155 978 -155 1 s2o
rlabel metal1 842 -1014 842 -1014 1 clk
rlabel metal1 911 -1010 911 -1010 1 clk
rlabel metal1 957 -1011 957 -1011 1 clk
rlabel metal1 979 -1010 979 -1010 1 clk
rlabel metal1 924 -826 924 -826 1 vdd
rlabel metal1 1016 -1082 1016 -1082 1 gnd
rlabel metal1 1045 -916 1045 -916 1 s4o
rlabel metal1 735 -1446 735 -1446 1 clk
rlabel metal1 804 -1442 804 -1442 1 clk
rlabel metal1 850 -1443 850 -1443 1 clk
rlabel metal1 872 -1442 872 -1442 1 clk
rlabel metal1 817 -1258 817 -1258 1 vdd
rlabel metal1 909 -1514 909 -1514 1 gnd
rlabel metal1 941 -1347 941 -1347 1 c4o
rlabel metal1 311 -1625 311 -1625 7 gnd
rlabel metal1 55 -1717 55 -1717 7 vdd
rlabel metal1 239 -1662 239 -1662 7 clk
rlabel metal1 240 -1684 240 -1684 7 clk
rlabel metal1 239 -1730 239 -1730 7 clk
rlabel metal1 243 -1799 243 -1799 7 clk
rlabel metal1 165 -1816 165 -1816 1 b4i
rlabel metal2 118 -1320 118 -1320 1 a4
rlabel metal1 60 -1581 60 -1581 1 gnd
rlabel metal1 -32 -1325 -32 -1325 1 vdd
rlabel metal1 23 -1509 23 -1509 1 clk
rlabel metal1 1 -1510 1 -1510 1 clk
rlabel metal1 -45 -1509 -45 -1509 1 clk
rlabel metal1 -114 -1513 -114 -1513 1 clk
rlabel metal1 -132 -1471 -132 -1471 3 a4i
rlabel metal1 75 -1259 75 -1259 7 clk
rlabel metal1 71 -1190 71 -1190 7 clk
rlabel metal1 72 -1144 72 -1144 7 clk
rlabel metal1 71 -1122 71 -1122 7 clk
rlabel metal1 -113 -1177 -113 -1177 7 vdd
rlabel metal1 143 -1085 143 -1085 7 gnd
rlabel metal1 32 -1278 34 -1276 1 b3i
rlabel metal1 -112 -903 -112 -903 1 clk
rlabel metal1 -43 -899 -43 -899 1 clk
rlabel metal1 3 -900 3 -900 1 clk
rlabel metal1 25 -899 25 -899 1 clk
rlabel metal1 -30 -715 -30 -715 1 vdd
rlabel metal1 62 -971 62 -971 1 gnd
rlabel metal1 -129 -850 -129 -850 1 a3i
rlabel metal1 1052 -488 1052 -488 1 s3o
rlabel metal1 1023 -654 1023 -654 1 gnd
rlabel metal1 931 -398 931 -398 1 vdd
rlabel metal1 986 -582 986 -582 1 clk
rlabel metal1 964 -583 964 -583 1 clk
rlabel metal1 918 -582 918 -582 1 clk
rlabel metal1 849 -586 849 -586 1 clk
rlabel metal1 42 -692 42 -692 1 gnd
rlabel metal1 -50 -436 -50 -436 1 vdd
rlabel metal1 5 -620 5 -620 1 clk
rlabel metal1 -17 -621 -17 -621 1 clk
rlabel metal1 -63 -620 -63 -620 1 clk
rlabel metal1 -132 -624 -132 -624 1 clk
rlabel metal1 -150 -618 -150 -618 3 b2i
rlabel metal1 -193 -380 -193 -380 3 gnd
rlabel metal1 63 -288 63 -288 3 vdd
rlabel metal1 -121 -343 -121 -343 3 clk
rlabel metal1 -122 -321 -122 -321 3 clk
rlabel metal1 -121 -275 -121 -275 3 clk
rlabel metal1 -125 -206 -125 -206 3 clk
rlabel metal1 306 57 306 57 3 gnd
rlabel metal1 562 149 562 149 3 vdd
rlabel metal1 378 94 378 94 3 clk
rlabel metal1 377 116 377 116 3 clk
rlabel metal1 378 162 378 162 3 clk
rlabel metal1 374 231 374 231 3 clk
rlabel metal1 473 25 473 25 1 c0
rlabel metal1 417 253 418 253 1 c0i
rlabel metal1 261 128 261 128 3 vdd
rlabel metal1 77 73 77 73 3 clk
rlabel metal1 76 95 76 95 3 clk
rlabel metal1 77 141 77 141 3 clk
rlabel metal1 73 210 73 210 3 clk
rlabel metal1 5 36 5 36 3 gnd
rlabel metal1 114 226 114 226 1 b1i
rlabel metal1 -40 -169 -40 -169 1 gnd
rlabel metal1 -214 -101 -214 -101 1 clk
rlabel metal1 -145 -97 -145 -97 1 clk
rlabel metal1 -99 -98 -99 -98 1 clk
rlabel metal1 -77 -97 -77 -97 1 clk
rlabel metal1 -132 87 -132 87 1 vdd
rlabel metal1 -230 -60 -230 -60 3 a1i
rlabel metal1 -74 -189 -74 -189 1 a2i
rlabel metal1 1050 -25 1050 -25 1 gnd
rlabel metal1 1061 228 1061 228 1 vdd
rlabel metal1 1061 -321 1061 -321 1 gnd
rlabel metal1 1072 -68 1072 -68 1 vdd
rlabel metal1 1128 -654 1128 -654 1 gnd
rlabel metal1 1139 -401 1139 -401 1 vdd
rlabel metal1 1128 -1082 1128 -1082 1 gnd
rlabel metal1 1139 -829 1139 -829 1 vdd
rlabel metal1 1021 -1514 1021 -1514 1 gnd
rlabel metal1 1032 -1261 1032 -1261 1 vdd
<< end >>

magic
tech scmos
timestamp 1731823769
<< nwell >>
rect 107 24 213 26
rect 237 24 307 26
rect 107 -34 307 24
rect 211 -36 242 -34
rect 103 -140 134 -80
rect 170 -134 201 -74
<< ntransistor >>
rect 227 -132 229 -112
rect 250 -131 252 -111
rect 267 -131 269 -111
rect 289 -131 291 -111
rect 116 -199 118 -179
rect 176 -199 178 -179
rect 221 -198 223 -178
rect 250 -198 252 -178
<< ptransistor >>
rect 120 -23 122 17
rect 172 -23 174 17
rect 224 -25 226 15
rect 250 -24 252 17
rect 267 -23 269 17
rect 289 -23 291 17
rect 116 -128 118 -89
rect 183 -122 185 -83
<< ndiffusion >>
rect 226 -132 227 -112
rect 229 -132 230 -112
rect 249 -131 250 -111
rect 252 -131 253 -111
rect 266 -131 267 -111
rect 269 -131 270 -111
rect 288 -131 289 -111
rect 291 -131 292 -111
rect 115 -199 116 -179
rect 118 -199 119 -179
rect 175 -199 176 -179
rect 178 -199 179 -179
rect 220 -198 221 -178
rect 223 -198 224 -178
rect 249 -198 250 -178
rect 252 -198 253 -178
<< pdiffusion >>
rect 119 -23 120 17
rect 122 -23 123 17
rect 171 -23 172 17
rect 174 -23 175 17
rect 223 -25 224 15
rect 226 -25 227 15
rect 249 -24 250 17
rect 252 -24 253 17
rect 266 -23 267 17
rect 269 -23 270 17
rect 288 -23 289 17
rect 291 -23 292 17
rect 115 -128 116 -89
rect 118 -128 119 -89
rect 182 -122 183 -83
rect 185 -122 186 -83
<< ndcontact >>
rect 222 -132 226 -112
rect 230 -132 234 -112
rect 245 -131 249 -111
rect 253 -131 257 -111
rect 262 -131 266 -111
rect 270 -131 274 -111
rect 284 -131 288 -111
rect 292 -131 296 -111
rect 111 -199 115 -179
rect 119 -199 123 -179
rect 171 -199 175 -179
rect 179 -199 183 -179
rect 216 -198 220 -178
rect 224 -198 228 -178
rect 245 -198 249 -178
rect 253 -198 257 -178
<< pdcontact >>
rect 115 -23 119 17
rect 123 -23 127 17
rect 167 -23 171 17
rect 175 -23 179 17
rect 219 -25 223 15
rect 227 -25 231 15
rect 245 -24 249 17
rect 253 -24 257 17
rect 262 -23 266 17
rect 270 -23 274 17
rect 284 -23 288 17
rect 292 -23 296 17
rect 111 -128 115 -89
rect 119 -128 123 -89
rect 178 -122 182 -83
rect 186 -122 190 -83
<< polysilicon >>
rect 120 17 122 20
rect 172 17 174 20
rect 224 15 226 18
rect 250 17 252 20
rect 267 17 269 20
rect 289 17 291 20
rect 120 -45 122 -23
rect 172 -67 174 -23
rect 164 -69 174 -67
rect 224 -68 226 -25
rect 116 -89 118 -86
rect 116 -156 118 -128
rect 164 -162 166 -69
rect 216 -70 226 -68
rect 183 -83 185 -80
rect 183 -152 185 -122
rect 216 -162 218 -70
rect 250 -94 252 -24
rect 238 -96 252 -94
rect 227 -112 229 -109
rect 227 -153 229 -132
rect 164 -164 178 -162
rect 216 -164 223 -162
rect 116 -179 118 -176
rect 176 -179 178 -164
rect 221 -178 223 -164
rect 238 -172 240 -96
rect 250 -111 252 -108
rect 267 -111 269 -23
rect 289 -111 291 -23
rect 250 -151 252 -131
rect 267 -135 269 -131
rect 289 -134 291 -131
rect 238 -174 252 -172
rect 250 -178 252 -174
rect 116 -213 118 -199
rect 176 -213 178 -199
rect 221 -211 223 -198
rect 250 -213 252 -198
<< polycontact >>
rect 116 -45 120 -41
rect 168 -43 172 -39
rect 220 -58 224 -54
rect 246 -58 250 -54
rect 112 -156 116 -152
rect 179 -152 183 -148
rect 263 -58 267 -54
rect 223 -153 227 -149
rect 285 -58 289 -54
rect 246 -151 250 -147
rect 112 -212 116 -208
<< metal1 >>
rect 100 24 307 42
rect 115 17 119 24
rect 167 17 171 24
rect 97 -45 116 -41
rect 123 -57 127 -23
rect 111 -61 127 -57
rect 158 -43 168 -39
rect 111 -89 115 -61
rect 119 -152 123 -128
rect 158 -152 162 -43
rect 175 -50 179 -23
rect 219 15 223 24
rect 245 17 249 24
rect 262 17 266 24
rect 284 17 288 24
rect 175 -56 182 -50
rect 227 -54 231 -25
rect 253 -54 257 -24
rect 270 -54 274 -23
rect 292 -54 296 -23
rect 178 -83 182 -56
rect 208 -58 220 -54
rect 227 -58 246 -54
rect 253 -58 263 -54
rect 270 -58 285 -54
rect 292 -58 368 -54
rect 186 -148 190 -122
rect 208 -148 212 -58
rect 227 -76 231 -58
rect 222 -80 231 -76
rect 222 -112 226 -80
rect 253 -100 257 -58
rect 270 -98 274 -58
rect 292 -60 300 -58
rect 245 -104 257 -100
rect 262 -102 274 -98
rect 296 -100 300 -60
rect 245 -111 249 -104
rect 262 -111 266 -102
rect 284 -104 300 -100
rect 284 -111 288 -104
rect 174 -152 179 -148
rect 186 -152 212 -148
rect 105 -156 112 -152
rect 119 -156 162 -152
rect 119 -170 123 -156
rect 186 -168 190 -152
rect 220 -153 223 -149
rect 111 -174 123 -170
rect 171 -172 190 -168
rect 230 -169 234 -132
rect 243 -151 246 -147
rect 253 -165 257 -131
rect 111 -179 115 -174
rect 171 -179 175 -172
rect 216 -173 234 -169
rect 245 -169 257 -165
rect 216 -178 220 -173
rect 245 -178 249 -169
rect 103 -212 112 -208
rect 119 -216 123 -199
rect 179 -216 183 -199
rect 224 -216 228 -198
rect 253 -216 257 -198
rect 270 -216 274 -131
rect 292 -216 296 -131
rect 110 -228 314 -216
<< metal2 >>
rect 223 -153 227 -149
rect 246 -151 250 -147
<< labels >>
rlabel metal1 112 -43 112 -43 1 d
rlabel metal1 116 31 116 31 1 vdd
rlabel metal1 108 -210 108 -210 1 d
rlabel metal1 107 -154 107 -154 1 clk
rlabel metal1 310 -57 310 -57 1 qf
rlabel metal1 244 -149 244 -149 1 clk
rlabel metal1 221 -151 221 -151 1 clk
rlabel metal1 176 -150 176 -150 1 clk
rlabel metal1 285 -218 285 -218 1 gnd
rlabel metal1 269 -223 269 -223 1 gnd
<< end >>

* prelayout
.include TSMC_180nm.txt

.param LAMBDA=0.09u
.param SUPPLY=1.8
.param width=1.8u
.param Wp = 2*width
.param Wn = width
.global gnd vdd

Vdd vdd gnd 'SUPPLY'
Va1 a1i gnd pulse(0 0 1n 0 0 1n 2n)
Va2 a2i gnd pulse(0 0 1n 0 0 2n 4n)
Va3 a3i gnd pulse(0 0 1n 0 0 4n 8n)
Va4 a4i gnd pulse(0 0 1n 0 0 8n 16n)

Vb4 b4i gnd pulse(1.8 1.8 1n 0 0 16n 32n)
Vb3 b3i gnd pulse(1.8 1.8 1n 0 0 32n 64n)
Vb2 b2i gnd pulse(1.8 1.8 1n 0 0 64n 128n)
Vb1 b1i gnd pulse(1.8 1.8 1n 0 0 128n 256n)

Vcin c0i gnd pulse(0 0 1n 0 0 1n 2n)

Vclk clk gnd pulse(0 1.8 0.2n 0 0 0.5n 1n)


* Vb1 b1i gnd pulse(0 1.8 2n 0 0 32n 64n)
* Vb2 b2i gnd pulse(0 1.8 2n 0 0 64n 128n)
* Vb3 b3i gnd pulse(0 1.8 2n 0 0 128n 256n)
* Vb4 b4i gnd pulse(0 1.8 2n 0 0 256n 512n) 

.subckt tspc q_out d clk vdd gnd
M1 c d vdd vdd CMOSP W={wp} L={2*LAMBDA} 
+AS={5*wp*LAMBDA} PS={10*LAMBDA+2*wp} 
+AD={5*wp*LAMBDA} PD={10*LAMBDA+2*wp}
M2 out clk c vdd CMOSP W={wp} L={2*LAMBDA} 
+AS={5*wp*LAMBDA} PS={10*LAMBDA+2*wp} 
+AD={5*wp*LAMBDA} PD={10*LAMBDA+2*wp}
M3 out d gnd gnd CMOSN W={wn} L={2*LAMBDA} 
+AS={5*wn*LAMBDA} PS={10*LAMBDA+2*wn} 
+AD={5*wn*LAMBDA} PD={10*LAMBDA+2*wn}
M4 k out vdd vdd CMOSP W={wp} L={2*LAMBDA} 
+AS={5*wp*LAMBDA} PS={10*LAMBDA+2*wp} 
+AD={5*wp*LAMBDA} PD={10*LAMBDA+2*wp}
M5 f clk k vdd CMOSP W={wp} L={2*LAMBDA} 
+AS={5*wp*LAMBDA} PS={10*LAMBDA+2*wp} 
+AD={5*wp*LAMBDA} PD={10*LAMBDA+2*wp}
M6 f out gnd gnd CMOSN W={wn} L={2*LAMBDA} 
+AS={5*wn*LAMBDA} PS={10*LAMBDA+2*wn} 
+AD={5*wn*LAMBDA} PD={10*LAMBDA+2*wn}
M7 g f vdd vdd CMOSP W={wp} L={2*LAMBDA} 
+AS={5*wp*LAMBDA} PS={10*LAMBDA+2*wp} 
+AD={5*wp*LAMBDA} PD={10*LAMBDA+2*wp}
M8 g clk h gnd CMOSN W={wn} L={2*LAMBDA} 
+AS={5*wn*LAMBDA} PS={10*LAMBDA+2*wn} 
+AD={5*wn*LAMBDA} PD={10*LAMBDA+2*wn}
M9 h f gnd gnd CMOSN W={wn} L={2*LAMBDA} 
+AS={5*wn*LAMBDA} PS={10*LAMBDA+2*wn} 
+AD={5*wn*LAMBDA} PD={10*LAMBDA+2*wn}
M10 q g vdd vdd CMOSP W={wp} L={2*LAMBDA} 
+AS={5*wp*LAMBDA} PS={10*LAMBDA+2*wp} 
+AD={5*wp*LAMBDA} PD={10*LAMBDA+2*wp}
M11  q clk in gnd CMOSN W={wn} L={2*LAMBDA} 
+AS={5*wn*LAMBDA} PS={10*LAMBDA+2*wn} 
+AD={5*wn*LAMBDA} PD={10*LAMBDA+2*wn}
M12 in g gnd gnd CMOSN W={wn} L={2*LAMBDA} 
+AS={5*wn*LAMBDA} PS={10*LAMBDA+2*wn} 
+AD={5*wn*LAMBDA} PD={10*LAMBDA+2*wn}
Xinv1 out_not q vdd gnd inv
Xinv2 q_out out_not vdd gnd inv
.ends 

.subckt and y_bar a b vdd gnd
M1 y a vdd vdd CMOSP W={Wp} L={2*LAMBDA} 
+AS={5*Wp*LAMBDA} PS={10*LAMBDA+2*Wp} 
+AD={5*Wp*LAMBDA} PD={10*LAMBDA+2*Wp}
M3 y b vdd vdd CMOSP W={Wp} L={2*LAMBDA} 
+AS={5*Wp*LAMBDA} PS={10*LAMBDA+2*Wp} 
+AD={5*Wp*LAMBDA} PD={10*LAMBDA+2*Wp}
M2 y a w gnd CMOSN W={Wp} L={2*LAMBDA} 
+AS={5*Wp*LAMBDA} PS={10*LAMBDA+2*Wp} 
+AD={5*Wp*LAMBDA} PD={10*LAMBDA+2*Wp}
M4 w b gnd gnd CMOSN W={Wp} L={2*LAMBDA} 
+AS={5*Wp*LAMBDA} PS={10*LAMBDA+2*Wp} 
+AD={5*Wp*LAMBDA} PD={10*LAMBDA+2*Wp}
X1 y_bar y vdd gnd inv
.ends

.subckt xor y a b vdd gnd
X1 b_bar b vdd gnd inv
M1 y b a vdd CMOSP W={Wp} L={2*LAMBDA} 
+AS={5*Wp*LAMBDA} PS={10*LAMBDA+2*Wp} 
+AD={5*Wp*LAMBDA} PD={10*LAMBDA+2*Wp}
M2 y b_bar a gnd CMOSN W={Wn} L={2*LAMBDA} 
+AS={5*Wn*LAMBDA} PS={10*LAMBDA+2*Wn} 
+AD={5*Wn*LAMBDA} PD={10*LAMBDA+2*Wn}
M3 y a b vdd CMOSP W={Wp} L={2*LAMBDA} 
+AS={5*Wp*LAMBDA} PS={10*LAMBDA+2*Wp} 
+AD={5*Wp*LAMBDA} PD={10*LAMBDA+2*Wp}
M4 y a b_bar gnd CMOSN W={Wn} L={2*LAMBDA} 
+AS={5*Wn*LAMBDA} PS={10*LAMBDA+2*Wn} 
+AD={5*Wn*LAMBDA} PD={10*LAMBDA+2*Wn}
.ends

.subckt inv y x vdd gnd 
M1 y x vdd vdd CMOSP W={Wp} L={2*LAMBDA} 
+AS={5*Wp*LAMBDA} PS={10*LAMBDA+2*Wp} 
+AD={5*Wp*LAMBDA} PD={10*LAMBDA+2*Wp}
M2 y x gnd gnd CMOSN W={Wn} L={2*LAMBDA} 
+AS={5*Wn*LAMBDA} PS={10*LAMBDA+2*Wn} 
+AD={5*Wn*LAMBDA} PD={10*LAMBDA+2*Wn}
.ends

.subckt C1block  c1 p1 g1 c0  
M1  t1 p1 vdd vdd CMOSP W={2*Wp} L={2*LAMBDA} 
+AS={5*2*Wp*LAMBDA} PS={10*LAMBDA+2*Wp*2} 
+AD={5*Wp*2*LAMBDA} PD={10*LAMBDA+2*Wp*2}
M2 t1 c0 vdd vdd CMOSP  W={2*Wp} L={2*LAMBDA} 
+AS={5*2*Wp*LAMBDA} PS={10*LAMBDA+2*Wp*2} 
+AD={5*Wp*2*LAMBDA} PD={10*LAMBDA+2*Wp*2}
M3 c1_bar g1 t1 vdd CMOSP W={2*Wp} L={2*LAMBDA} 
+AS={5*2*Wp*LAMBDA} PS={10*LAMBDA+2*Wp*2} 
+AD={5*Wp*2*LAMBDA} PD={10*LAMBDA+2*Wp*2}

M4 c1_bar p1 t2 gnd CMOSN W={2*Wn} L={2*LAMBDA} 
+AS={5*2*Wn*LAMBDA} PS={10*LAMBDA+2*2*Wn} 
+AD={5*2*Wn*LAMBDA} PD={10*LAMBDA+2*2*Wn} 
M5 t2 c0 gnd gnd CMOSN W={2*Wn} L={2*LAMBDA} 
+AS={5*2*Wn*LAMBDA} PS={10*LAMBDA+2*2*Wn} 
+AD={5*2*Wn*LAMBDA} PD={10*LAMBDA+2*2*Wn} 
M6 c1_bar g1 gnd gnd CMOSN W={Wn} L={2*LAMBDA} 
+AS={5*Wn*LAMBDA} PS={10*LAMBDA+2*Wn} 
+AD={5*Wn*LAMBDA} PD={10*LAMBDA+2*Wn}
X1 c1 c1_bar vdd gnd inv

.ends

.subckt c2block p2 p1 g2 g1 c0 c2 
M1 t2 p2 vdd vdd CMOSP W={1.5*Wp} L={2*LAMBDA} 
+AS={5*1.5*Wp*LAMBDA} PS={10*LAMBDA+2*Wp*1.5} 
+AD={5*Wp*1.5*LAMBDA} PD={10*LAMBDA+2*Wp*1.5}
M2 c2_bar g2 t2 vdd CMOSP W={Wp*3} L={2*LAMBDA} 
+AS={5*Wp*3*LAMBDA} PS={10*LAMBDA+2*Wp*3} 
+AD={5*Wp*3*LAMBDA} PD={10*LAMBDA+2*Wp*3}
M3 t2 g1 t1 vdd CMOSP W={Wp*3} L={2*LAMBDA} 
+AS={5*Wp*3*LAMBDA} PS={10*LAMBDA+2*Wp*3} 
+AD={5*Wp*3*LAMBDA} PD={10*LAMBDA+2*Wp*3}
M4 t1 p1 vdd vdd CMOSP W={Wp*3} L={2*LAMBDA} 
+AS={5*Wp*3*LAMBDA} PS={10*LAMBDA+2*Wp*3} 
+AD={5*Wp*3*LAMBDA} PD={10*LAMBDA+2*Wp*3} 
M5 t1 c0 vdd vdd CMOSP W={Wp*3} L={2*LAMBDA} 
+AS={5*Wp*3*LAMBDA} PS={10*LAMBDA+2*Wp*3} 
+AD={5*Wp*3*LAMBDA} PD={10*LAMBDA+2*Wp*3}

M6 c2_bar p2 t3 gnd CMOSN W={3*Wn} L={2*LAMBDA} 
+AS={5*Wn*3*LAMBDA} PS={10*LAMBDA+2*Wn*3} 
+AD={5*Wn*3*LAMBDA} PD={10*LAMBDA+2*Wn*3}
M7 t3 p1 t4 gnd CMOSN W={3*Wn} L={2*LAMBDA} 
+AS={5*Wn*3*LAMBDA} PS={10*LAMBDA+2*Wn*3} 
+AD={5*Wn*3*LAMBDA} PD={10*LAMBDA+2*Wn*3}
M8 t4 c0 gnd gnd CMOSN W={3*Wn} L={2*LAMBDA} 
+AS={5*Wn*3*LAMBDA} PS={10*LAMBDA+2*Wn*3} 
+AD={5*Wn*3*LAMBDA} PD={10*LAMBDA+2*Wn*3}
M9 t3 g1 gnd gnd CMOSN W={1.5*Wn} L={2*LAMBDA} 
+AS={5*Wn*1.5*LAMBDA} PS={10*LAMBDA+2*Wn*1.5} 
+AD={5*Wn*1.5*LAMBDA} PD={10*LAMBDA+2*Wn*1.5}
M10 c2_bar g2 gnd gnd CMOSN W={Wn} L={2*LAMBDA} 
+AS={5*Wn*LAMBDA} PS={10*LAMBDA+2*Wn} 
+AD={5*Wn*LAMBDA} PD={10*LAMBDA+2*Wn}

X1 c2 c2_bar vdd gnd inv
.ends

.subckt c3block p3 p2 p1 g3 g2 g1 c0 c3 
M1 t3 p3 vdd vdd CMOSP W={Wp*1.33} L={2*LAMBDA} 
+AS={5*Wp*1.33*LAMBDA} PS={10*LAMBDA+2*Wp*1.33} 
+AD={5*Wp*1.33*LAMBDA} PD={10*LAMBDA+2*Wp*1.33}
M2 c3_bar g3 t3 vdd CMOSP W={Wp*4} L={2*LAMBDA} 
+AS={5*Wp*4*LAMBDA} PS={10*LAMBDA+2*Wp*4} 
+AD={5*Wp*4*LAMBDA} PD={10*LAMBDA+2*Wp*4}
M3 t2 p2 vdd vdd CMOSP  W={Wp*2} L={2*LAMBDA} 
+AS={5*Wp*2*LAMBDA} PS={10*LAMBDA+2*Wp*2} 
+AD={5*Wp*2*LAMBDA} PD={10*LAMBDA+2*Wp*2}
M4 t3 g2 t2 vdd CMOSP W={Wp*4} L={2*LAMBDA} 
+AS={5*Wp*4*LAMBDA} PS={10*LAMBDA+2*Wp*4} 
+AD={5*Wp*4*LAMBDA} PD={10*LAMBDA+2*Wp*4}
M5 t1 p1 vdd vdd CMOSP W={Wp*4} L={2*LAMBDA} 
+AS={5*Wp*4*LAMBDA} PS={10*LAMBDA+2*Wp*4} 
+AD={5*Wp*4*LAMBDA} PD={10*LAMBDA+2*Wp*4}
M6 t1 c0 vdd vdd CMOSP W={Wp*4} L={2*LAMBDA} 
+AS={5*Wp*4*LAMBDA} PS={10*LAMBDA+2*Wp*4} 
+AD={5*Wp*4*LAMBDA} PD={10*LAMBDA+2*Wp*4}
M7 t2 g1 vdd vdd CMOSP W={Wp*4} L={2*LAMBDA} 
+AS={5*Wp*4*LAMBDA} PS={10*LAMBDA+2*Wp*4} 
+AD={5*Wp*4*LAMBDA} PD={10*LAMBDA+2*Wp*4}


M8 c3_bar p3 t4 gnd CMOSN W={4*Wn} L={2*LAMBDA} 
+AS={5*Wn*4*LAMBDA} PS={10*LAMBDA+2*Wn*4} 
+AD={5*Wn*4*LAMBDA} PD={10*LAMBDA+2*Wn*4}
M9 t4 p2 t5 gnd CMOSN W={4*Wn} L={2*LAMBDA} 
+AS={5*Wn*4*LAMBDA} PS={10*LAMBDA+2*Wn*4} 
+AD={5*Wn*4*LAMBDA} PD={10*LAMBDA+2*Wn*4}
M10 t5 p1 t6 gnd CMOSN W={4*Wn} L={2*LAMBDA} 
+AS={5*Wn*4*LAMBDA} PS={10*LAMBDA+2*Wn*4} 
+AD={5*Wn*4*LAMBDA} PD={10*LAMBDA+2*Wn*4}
M11 t6 c0 gnd gnd CMOSN W={4*Wn} L={2*LAMBDA} 
+AS={5*Wn*4*LAMBDA} PS={10*LAMBDA+2*Wn*4} 
+AD={5*Wn*4*LAMBDA} PD={10*LAMBDA+2*Wn*4}
M12 t5 g1 gnd gnd CMOSN W={2*Wn} L={2*LAMBDA} 
+AS={5*Wn*2*LAMBDA} PS={10*LAMBDA+2*2*Wn} 
+AD={5*Wn*2*LAMBDA} PD={10*LAMBDA+2*Wn*2}
M13 t4 g2 gnd gnd CMOSN W={1.33*Wn} L={2*LAMBDA} 
+AS={5*Wn*1.33*LAMBDA} PS={10*LAMBDA+2*Wn*1.33} 
+AD={5*Wn*1.33*LAMBDA} PD={10*LAMBDA+2*Wn*1.33}
M14 c3_bar g3 gnd gnd CMOSN W={Wn} L={2*LAMBDA} 
+AS={5*Wn*LAMBDA} PS={10*LAMBDA+2*Wn} 
+AD={5*Wn*LAMBDA} PD={10*LAMBDA+2*Wn}

X1 c3 c3_bar vdd gnd inv
.ends

.subckt c4block p4 p3 p2 p1 g4 g3 g2 g1 c0 c4
M1 t4 p4 vdd vdd CMOSP W={Wp*1.25} L={2*LAMBDA} 
+AS={5*Wp*1.25*LAMBDA} PS={10*LAMBDA+2*Wp*1.25} 
+AD={5*Wp*1.25*LAMBDA} PD={10*LAMBDA+2*Wp*1.25}
M2 c4_bar g4 t4 vdd CMOSP W={Wp*5} L={2*LAMBDA} 
+AS={5*Wp*5*LAMBDA} PS={10*LAMBDA+2*Wp*5} 
+AD={5*Wp*5*LAMBDA} PD={10*LAMBDA+2*Wp*5}
M3 t3 p3 vdd vdd CMOSP W={Wp*1.66} L={2*LAMBDA} 
+AS={5*Wp*1.66*LAMBDA} PS={10*LAMBDA+2*Wp*1.66} 
+AD={5*Wp*1.66*LAMBDA} PD={10*LAMBDA+2*Wp*1.66} 
M4 t4 g3 t3 vdd CMOSP W={Wp*5} L={2*LAMBDA} 
+AS={5*Wp*5*LAMBDA} PS={10*LAMBDA+2*Wp*5} 
+AD={5*Wp*5*LAMBDA} PD={10*LAMBDA+2*Wp*5}
M5 t2 p2 vdd vdd CMOSP W={Wp*2.5} L={2*LAMBDA} 
+AS={5*Wp*2.5*LAMBDA} PS={10*LAMBDA+2*Wp*2.5} 
+AD={5*Wp*2.5*LAMBDA} PD={10*LAMBDA+2*Wp*2.5}
M6 t3 g2 t2 vdd CMOSP W={Wp*5} L={2*LAMBDA} 
+AS={5*Wp*5*LAMBDA} PS={10*LAMBDA+2*Wp*5} 
+AD={5*Wp*5*LAMBDA} PD={10*LAMBDA+2*Wp*5}
M7 t1 p1 vdd vdd CMOSP W={Wp*5} L={2*LAMBDA} 
+AS={5*Wp*5*LAMBDA} PS={10*LAMBDA+2*Wp*5} 
+AD={5*Wp*5*LAMBDA} PD={10*LAMBDA+2*Wp*5}
M8 t2 g1 t1 vdd CMOSP W={Wp*5} L={2*LAMBDA} 
+AS={5*Wp*5*LAMBDA} PS={10*LAMBDA+2*Wp*5} 
+AD={5*Wp*5*LAMBDA} PD={10*LAMBDA+2*Wp*5} 
M9 t1 c0 vdd vdd CMOSP W={Wp*5} L={2*LAMBDA} 
+AS={5*Wp*5*LAMBDA} PS={10*LAMBDA+2*Wp*5} 
+AD={5*Wp*5*LAMBDA} PD={10*LAMBDA+2*Wp*5}

M10 c4_bar p4 t5 gnd CMOSN  W={Wn*5} L={2*LAMBDA} 
+AS={5*Wn*5*LAMBDA} PS={10*LAMBDA+2*Wn*5} 
+AD={5*Wn*5*LAMBDA} PD={10*LAMBDA+2*Wn*5}
M11 t5 p3 t6 gnd CMOSN W={Wn*5} L={2*LAMBDA} 
+AS={5*Wn*5*LAMBDA} PS={10*LAMBDA+2*Wn*5} 
+AD={5*Wn*5*LAMBDA} PD={10*LAMBDA+2*Wn*5}
M12 t6 p2 t7 gnd CMOSN W={Wn*5} L={2*LAMBDA} 
+AS={5*Wn*5*LAMBDA} PS={10*LAMBDA+2*Wn*5} 
+AD={5*Wn*5*LAMBDA} PD={10*LAMBDA+2*Wn*5}
M13 t7 p1 t8 gnd CMOSN W={Wn*5} L={2*LAMBDA} 
+AS={5*Wn*5*LAMBDA} PS={10*LAMBDA+2*Wn*5} 
+AD={5*Wn*5*LAMBDA} PD={10*LAMBDA+2*Wn*5}
M14 t8 c0 gnd gnd CMOSN W={Wn*5} L={2*LAMBDA} 
+AS={5*Wn*5*LAMBDA} PS={10*LAMBDA+2*Wn*5} 
+AD={5*Wn*5*LAMBDA} PD={10*LAMBDA+2*Wn*5}
M15 t7 g1 gnd gnd CMOSN W={Wn*2.5} L={2*LAMBDA} 
+AS={5*Wn*2.5*LAMBDA} PS={10*LAMBDA+2*Wn*2.5} 
+AD={5*Wn*2.5*LAMBDA} PD={10*LAMBDA+2*Wn*2.5}
M16 t6 g2 gnd gnd CMOSN W={Wn*1.66} L={2*LAMBDA} 
+AS={5*Wn*1.66*LAMBDA} PS={10*LAMBDA+2*Wn*1.66} 
+AD={5*Wn*1.66*LAMBDA} PD={10*LAMBDA+2*Wn*1.66}
M17 t5 g3 gnd gnd CMOSN W={Wn*1.25} L={2*LAMBDA} 
+AS={5*Wn*1.25*LAMBDA} PS={10*LAMBDA+2*Wn*1.25} 
+AD={5*Wn*1.25*LAMBDA} PD={10*LAMBDA+2*Wn*1.25}
M18 c4_bar g4 gnd gnd CMOSN W={Wn} L={2*LAMBDA} 
+AS={5*Wn*LAMBDA} PS={10*LAMBDA+2*Wn} 
+AD={5*Wn*LAMBDA} PD={10*LAMBDA+2*Wn}

X1 c4 c4_bar vdd gnd inv
.ends


x17 a1 a1i clk vdd gnd tspc 
x18 a2 a2i clk vdd gnd tspc
x19 a3 a3i clk vdd gnd tspc
x20 a4 a4i clk vdd gnd tspc

x21 b1 b1i clk vdd gnd tspc
x22 b2 b2i clk vdd gnd tspc
x23 b3 b3i clk vdd gnd tspc
x24 b4 b4i clk vdd gnd tspc
x25 c0 c0i clk vdd gnd tspc
* propogates
X1 p1 a1 b1 vdd gnd xor
X2 p2 a2 b2 vdd gnd xor
X3 p3 a3 b3 vdd gnd xor
X4 p4 a4 b4 vdd gnd xor

* * * generates
X5 g1 a1 b1 vdd gnd and
X6 g2 a2 b2 vdd gnd and
X7 g3 a3 b3 vdd gnd and
X8 g4 a4 b4 vdd gnd and

* carry
X9  c1 p1 g1 c0 c1block
X10 p2 p1 g2 g1 c0 c2 C2block
X11 p3 p2 p1 g3 g2 g1 c0 c3 c3block
X12 p4 p3 p2 p1 g4 g3 g2 g1 c0 c4 c4block

* sum
X13 s1 p1 c0 vdd gnd xor
X14 s2 p2 c1 vdd gnd xor
X15 s3 p3 c2 vdd gnd xor
X16 s4 p4 c3 vdd gnd xor

x26 s1o s1 clk vdd gnd tspc
x27 s2o s2 clk vdd gnd tspc
x28 s3o s3 clk vdd gnd tspc
x29 s4o s4 clk vdd gnd tspc
x35 c4o c4 clk vdd gnd tspc
* inverters in the end
x30 y1 c4 vdd gnd inv
x31 y2 s4 vdd gnd inv 
x32 y3 s3 vdd gnd inv
x33 y4 s2 vdd gnd inv
x34 y5 s1 vdd gnd inv
.measure tran delays0 TRIG v(c0) VAL=0.9 RISE=1 TARG v(c4) VAL=0.9 rise=1
.tran 0.1n 50n

.control
set hcopypscolor=1
set color0=white
set color1=black
run
set curplottitle="Sanjana Sheela - 20231012027- prelayout"
* plot v(a1i) v(a2i)+2 v(a3i)+4 v(a4i)+6 v(clk)+8
* plot v(b1i) v(b2i)+2 v(b3i)+4 v(b4i)+6 v(clk)+8 v(c0i)-2
* plot v(a1) v(a2)+2 v(a3)+4 v(a4)+6 v(clk)+8 v(c0)-2
* plot v(b1) v(b2)+2 v(b3)+4 v(b4)+6 v(clk)+8 v(c0)-2
plot v(s1o) v(s2o)+2 v(s3o)+4 v(s4o)+6 v(c4o)+8 v(clk)+10
* plot v(g1) v(p1)+2 v(g2)+4 v(p2)+6 v(g3)+8 v(p3)+10 v(g4)+12 v(p4)+14
* plot v(c0)-2 v(c1) v(c2)+2 v(c3)+4 v(c4)+6
* plot v(s1) v(s2)+2 v(s3)+4 v(s4)+6 v(c4)+8

* plot v(a1i) v(a1)+2 v(clk)+4
* plot v(a2i) v(a2)+2 v(clk)+4
* plot v(a3i) v(a3)+2 v(clk)+4
* plot v(a4i) v(a4)+2 v(clk)+4

* plot v(b1i) v(b1)+2 v(clk)+4
* plot v(b2i) v(b2)+2 v(clk)+4
* plot v(b3i) v(b3)+2 v(clk)+4
* plot v(b4i) v(b4)+2 v(clk)+4

* plot v(c0i) v(c0)+2 v(clk)+4

* plot v(s1) v(s1o)+2 v(clk)+4
* plot v(s2) v(s2o)+2 v(clk)+4
* plot v(s3) v(s3o)+2 v(clk)+4
* plot v(s4) v(s4o)+2 v(clk)+4

* plot v(a1) v(b1)+2 v(p1)+4 
* plot v(a2) v(b2)+2 v(p2)+4 
* plot v(a3) v(b3)+2 v(p3)+4 
* plot v(a4) v(b4)+2 v(p4)+4

* plot v(a1) v(b1)+2 v(g1)+4 
* plot v(a2) v(b2)+2 v(g2)+4 
* plot v(a3) v(b3)+2 v(g3)+4 
* plot v(a4) v(b4)+2 v(g4)+4

* plot v(p1) v(g1)+2 v(c0)+4 v(c1)+6
* plot v(p2) v(g2)+2 v(c1)+4 v(c2)+6
* plot v(p3) v(g3)+2 v(c2)+4 v(c3)+6
* plot v(p4) v(g4)+2 v(c3)+4 v(c4)+6
* plot v(c2) v(p3)+2 v(s3)+4

* plot v(a1) v(b1)+2 v(c0)+4 v(p1)+6 v(g1)+8 v(s1)+10 v(c1)+12
* plot v(a2) v(b2)+2 v(c1)+4 v(p2)+6 v(g2)+8 v(s2)+10 v(c2)+12
* plot v(a3) v(b3)+2 v(c2)+4 v(p3)+6 v(g3)+8 v(s3)+10 v(c3)+12
* plot v(a4) v(b4)+2 v(c3)+4 v(p4)+6 v(g4)+8 v(s4)+10 v(c4)+12

.endc
.end

* 
.include TSMC_180nm.txt

.param LAMBDA=0.09u
.param SUPPLY=1.8
.param width=1.8u
.param Wp = 2*width
.param Wn = width
.global gnd vdd

VD1 vdd1 0 1.8V
VD2 vdd11 0 1.8V
VD3 vdd2 0 1.8V
VD4 vdd22 0 1.8V
VD5 vddc1 0 1.8V
VD6 vddc2 0 1.8V
VD7 vdd33 0 1.8V
VD8 vdd3 0 1.8V
VD9 vddc3 0 1.8V
VD10 vdd44 0 1.8V
VD11 vdd4 0 1.8V
VD12 vddc4 0 1.8V

VG1 gnd1 0 0
VG2 gnd11 0 0
VG3 gnd2 0 0
VG4 gnd22 0 0
VG5 gndc2 0 0
VG6 gndc1 0 0
VG7 gnd3 0 0
VG8 gnd33 0 0
VG9 gndc3 0 0
VG10 gnd4 0 0
VG11 gnd44 0 0
VG12 gndc4 0 0

Vdd vdd gnd 'SUPPLY'
Va1 p1 gnd pulse(0 1.8 2n 0 0 2n 4n)
Va2 p2 gnd pulse(0 1.8 2n 0 0 4n 8n)
Va3 p3 gnd pulse(0 1.8 2n 0 0 8n 16n)
Va4 p4 gnd pulse(0 1.8 2n 0 0 16n 32n)

Vb1 g1 gnd pulse(0 1.8 2n 0 0 16n 32n)
Vb2 g2 gnd pulse(0 1.8 2n 0 0 8n 16n)
Vb3 g3 gnd pulse(0 1.8 2n 0 0 4n 8n)
Vb4 g4 gnd pulse(0 1.8 2n 0 0 2n 4n)
Vin c0 gnd pulse(0 1.8 2n 0 0 2n 4n)

* SPICE3 file created from carryblock.ext - technology: scmos

.option scale=0.09u

M1000 gndc1 g1 a_681_n251# Gnd CMOSN w=20 l=2
+  ad=400 pd=190 as=300 ps=140
M1001 gndc3 g1 a_579_n1432# Gnd CMOSN w=40 l=2
+  ad=930 pd=422 as=1000 ps=430
M1002 c2 a_688_n831# vddc2 w_626_n700# CMOSP w=40 l=2
+  ad=200 pd=90 as=1700 ps=720
M1003 a_634_n1180# GG a_597_n1181# w_545_n1187# CMOSP w=160 l=2
+  ad=1870 pd=778 as=2000 ps=830
M1004 vddc4 p3 a_623_n1911# w_538_n1918# CMOSP w=66 l=2
+  ad=3280 pd=1372 as=2330 ps=962
M1005 c4 a_678_n2188# gndc4 Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=1240 ps=556
M1006 vddc2 p1 a_639_n692# w_626_n700# CMOSP w=120 l=2
+  ad=0 pd=0 as=1800 ps=510
M1007 a_551_n2188# c0 gndc4 Gnd CMOSN w=100 l=2
+  ad=1000 pd=420 as=0 ps=0
M1008 a_678_n2188# g4 a_659_n1911# w_538_n1918# CMOSP w=200 l=2
+  ad=1000 pd=410 as=2250 ps=930
M1009 a_570_n2188# p1 a_551_n2188# Gnd CMOSN w=100 l=2
+  ad=1250 pd=530 as=0 ps=0
M1010 a_641_n2188# p3 a_606_n2188# Gnd CMOSN w=100 l=2
+  ad=1125 pd=480 as=1165 ps=496
M1011 vddc4 p2 a_588_n1911# w_538_n1918# CMOSP w=100 l=2
+  ad=0 pd=0 as=2500 ps=1030
M1012 gndc4 GG a_606_n2188# Gnd CMOSN w=33 l=2
+  ad=0 pd=0 as=0 ps=0
M1013 gndc2 g1 a_651_n831# Gnd CMOSN w=30 l=2
+  ad=650 pd=300 as=750 ps=330
M1014 a_597_n1181# g1 a_561_n1181# w_545_n1187# CMOSP w=160 l=2
+  ad=0 pd=0 as=2400 ps=990
M1015 gndc3 GG a_615_n1432# Gnd CMOSN w=26 l=2
+  ad=0 pd=0 as=930 ps=402
M1016 gndc3 g3 a_653_n1431# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=500 ps=220
M1017 a_653_n1431# p3 a_615_n1432# Gnd CMOSN w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1018 c1 a_681_n251# gndc1 Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1019 a_639_n831# c0 gndc2 Gnd CMOSN w=60 l=2
+  ad=600 pd=140 as=0 ps=0
M1020 a_681_n251# p1 a_664_n251# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1021 a_653_n1431# g3 a_634_n1180# w_545_n1187# CMOSP w=160 l=2
+  ad=800 pd=330 as=0 ps=0
M1022 c1 a_681_n251# vddc1 w_644_n126# CMOSP w=40 l=2
+  ad=200 pd=90 as=1000 ps=430
M1023 a_561_n1431# c0 gndc3 Gnd CMOSN w=80 l=2
+  ad=800 pd=340 as=0 ps=0
M1024 a_579_n1432# p1 a_561_n1431# Gnd CMOSN w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1025 a_688_n831# p2 a_651_n831# Gnd CMOSN w=60 l=2
+  ad=400 pd=180 as=0 ps=0
M1026 gndc4 g1 a_570_n2188# Gnd CMOSN w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 gndc4 a_652_n2046# a_641_n2188# Gnd CMOSN w=25 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 a_651_n831# p1 a_639_n831# Gnd CMOSN w=60 l=2
+  ad=0 pd=0 as=0 ps=0
M1029 c3 a_653_n1431# gndc3 Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1030 a_678_n2188# p4 a_641_n2188# Gnd CMOSN w=100 l=2
+  ad=600 pd=260 as=0 ps=0
M1031 vddc1 p1 a_664_n120# w_644_n126# CMOSP w=80 l=2
+  ad=0 pd=0 as=1200 ps=510
M1032 vddc2 p2 a_670_n693# w_626_n700# CMOSP w=60 l=2
+  ad=0 pd=0 as=1500 ps=630
M1033 vddc4 p4 a_659_n1911# w_538_n1918# CMOSP w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 gndc4 g4 a_678_n2188# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1035 a_551_n1911# c0 vddc4 w_538_n1918# CMOSP w=200 l=2
+  ad=3000 pd=1230 as=0 ps=0
M1036 a_681_n251# g1 a_664_n120# w_644_n126# CMOSP w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1037 a_670_n693# g1 a_639_n692# w_626_n700# CMOSP w=120 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 a_561_n1181# c0 vddc3 w_545_n1187# CMOSP w=160 l=2
+  ad=0 pd=0 as=2470 ps=1038
M1039 a_606_n2188# p2 a_570_n2188# Gnd CMOSN w=100 l=2
+  ad=0 pd=0 as=0 ps=0
M1040 vddc4 p1 a_551_n1911# w_538_n1918# CMOSP w=200 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 a_664_n251# c0 gndc1 Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1042 a_623_n1911# GG a_588_n1911# w_538_n1918# CMOSP w=200 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 gndc2 GG a_688_n831# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 a_688_n831# GG a_670_n693# w_626_n700# CMOSP w=120 l=2
+  ad=600 pd=250 as=0 ps=0
M1045 a_615_n1432# p2 a_579_n1432# Gnd CMOSN w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 a_664_n120# c0 vddc1 w_644_n126# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1047 vddc3 p2 a_597_n1181# w_545_n1187# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 c4 a_678_n2188# vddc4 w_538_n1918# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1049 a_639_n692# c0 vddc2 w_626_n700# CMOSP w=120 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 vddc3 p1 a_561_n1181# w_545_n1187# CMOSP w=160 l=2
+  ad=0 pd=0 as=0 ps=0
M1051 c3 a_653_n1431# vddc3 w_545_n1187# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1052 c2 a_688_n831# gndc2 Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1053 vddc3 p3 a_634_n1180# w_545_n1187# CMOSP w=54 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 a_588_n1911# g1 a_551_n1911# w_538_n1918# CMOSP w=200 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 a_659_n1911# a_652_n2046# a_623_n1911# w_538_n1918# CMOSP w=200 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_626_n700# vddc2 0.75fF
C1 g3 c0 0.20fF
C2 p4 w_538_n1918# 0.94fF
C3 vddc4 a_623_n1911# 1.13fF
C4 p2 g4 0.09fF
C5 GG g3 0.18fF
C6 p3 g3 0.18fF
C7 p2 g1 0.42fF
C8 a_651_n831# g1 0.08fF
C9 w_545_n1187# c3 0.46fF
C10 p2 p1 0.42fF
C11 GG c0 0.42fF
C12 gndc4 a_606_n2188# 0.71fF
C13 c1 gndc1 0.21fF
C14 p3 c0 0.29fF
C15 a_659_n1911# w_538_n1918# 0.56fF
C16 w_545_n1187# vddc3 0.92fF
C17 vddc2 c2 0.41fF
C18 p2 a_670_n693# 0.08fF
C19 vddc4 a_551_n1911# 5.55fF
C20 c2 gndc2 0.24fF
C21 GG p3 0.29fF
C22 w_545_n1187# g1 0.06fF
C23 GG a_606_n2188# 0.08fF
C24 gndc3 a_653_n1431# 0.21fF
C25 w_545_n1187# p1 0.06fF
C26 a_623_n1911# a_659_n1911# 2.06fF
C27 vddc3 a_597_n1181# 1.44fF
C28 a_678_n2188# g4 0.13fF
C29 w_626_n700# a_688_n831# 0.35fF
C30 w_644_n126# a_681_n251# 0.24fF
C31 a_615_n1432# a_653_n1431# 0.82fF
C32 w_538_n1918# c0 0.07fF
C33 w_545_n1187# a_653_n1431# 0.96fF
C34 vddc3 a_634_n1180# 1.07fF
C35 w_644_n126# g1 0.06fF
C36 GG w_538_n1918# 0.07fF
C37 p3 w_538_n1918# 0.85fF
C38 w_644_n126# p1 0.06fF
C39 a_681_n251# c1 0.07fF
C40 g4 a_652_n2046# 0.09fF
C41 vddc2 a_670_n693# 1.08fF
C42 gndc3 a_615_n1432# 0.42fF
C43 p3 a_623_n1911# 0.08fF
C44 a_688_n831# c2 0.08fF
C45 a_652_n2046# g1 0.09fF
C46 w_626_n700# c0 0.08fF
C47 a_652_n2046# p1 0.09fF
C48 vddc3 a_561_n1181# 4.50fF
C49 p4 g4 0.09fF
C50 a_588_n1911# w_538_n1918# 0.62fF
C51 a_634_n1180# a_653_n1431# 1.82fF
C52 w_545_n1187# p2 0.53fF
C53 w_626_n700# GG 0.07fF
C54 w_644_n126# vddc1 0.44fF
C55 a_561_n1181# p1 0.08fF
C56 p4 g1 0.09fF
C57 p4 p1 0.09fF
C58 gndc4 a_570_n2188# 1.01fF
C59 a_588_n1911# a_623_n1911# 2.06fF
C60 a_579_n1432# g1 0.08fF
C61 a_623_n1911# w_538_n1918# 0.57fF
C62 p2 a_597_n1181# 0.08fF
C63 a_678_n2188# c4 0.08fF
C64 vddc1 c1 0.41fF
C65 a_664_n120# a_681_n251# 0.91fF
C66 a_570_n2188# a_606_n2188# 1.03fF
C67 a_670_n693# a_688_n831# 1.24fF
C68 gndc2 a_651_n831# 0.78fF
C69 w_545_n1187# a_597_n1181# 0.50fF
C70 a_551_n1911# a_588_n1911# 2.13fF
C71 a_551_n1911# w_538_n1918# 0.71fF
C72 p1 a_664_n120# 0.09fF
C73 g3 g1 0.18fF
C74 g4 c0 0.09fF
C75 w_626_n700# a_639_n692# 0.21fF
C76 g3 p1 0.18fF
C77 p2 a_652_n2046# 0.09fF
C78 w_545_n1187# a_634_n1180# 0.54fF
C79 c4 vddc4 0.41fF
C80 gndc4 a_551_n2188# 1.26fF
C81 c0 g1 0.56fF
C82 GG g4 0.09fF
C83 p3 g4 0.09fF
C84 c0 p1 0.58fF
C85 p2 p4 0.09fF
C86 GG g1 0.42fF
C87 p3 g1 0.29fF
C88 gndc3 a_579_n1432# 0.70fF
C89 a_597_n1181# a_634_n1180# 1.65fF
C90 vddc1 a_664_n120# 1.80fF
C91 GG p1 0.42fF
C92 p3 p1 0.29fF
C93 g3 a_653_n1431# 0.17fF
C94 w_545_n1187# a_561_n1181# 0.55fF
C95 a_688_n831# a_651_n831# 0.62fF
C96 a_579_n1432# a_615_n1432# 0.82fF
C97 a_678_n2188# a_641_n2188# 1.03fF
C98 g4 w_538_n1918# 0.07fF
C99 a_561_n1181# a_597_n1181# 1.65fF
C100 w_538_n1918# g1 0.08fF
C101 w_626_n700# c2 0.08fF
C102 w_644_n126# c1 0.10fF
C103 a_664_n251# gndc1 0.41fF
C104 w_538_n1918# p1 0.08fF
C105 p2 g3 0.18fF
C106 gndc3 a_561_n1431# 0.82fF
C107 c4 gndc4 0.24fF
C108 a_641_n2188# a_652_n2046# 0.08fF
C109 a_639_n692# p1 0.06fF
C110 p2 c0 0.42fF
C111 a_681_n251# gndc1 0.24fF
C112 w_545_n1187# g3 0.08fF
C113 a_639_n692# a_670_n693# 1.24fF
C114 vddc2 a_688_n831# 0.02fF
C115 p2 GG 2.66fF
C116 a_678_n2188# a_659_n1911# 2.06fF
C117 a_688_n831# gndc2 0.26fF
C118 GG a_651_n831# 0.23fF
C119 p2 p3 0.29fF
C120 w_626_n700# g1 0.08fF
C121 p4 a_652_n2046# 0.09fF
C122 g1 gndc1 0.05fF
C123 w_545_n1187# c0 0.06fF
C124 w_626_n700# p1 0.08fF
C125 GG a_615_n1432# 0.08fF
C126 a_551_n1911# p1 0.08fF
C127 w_626_n700# a_670_n693# 0.42fF
C128 w_545_n1187# GG 0.07fF
C129 w_644_n126# a_664_n120# 0.35fF
C130 a_664_n251# a_681_n251# 0.41fF
C131 w_545_n1187# p3 0.69fF
C132 a_570_n2188# g1 0.09fF
C133 a_678_n2188# gndc4 0.33fF
C134 a_551_n2188# a_570_n2188# 1.03fF
C135 p2 a_588_n1911# 0.09fF
C136 c4 w_538_n1918# 0.54fF
C137 p2 w_538_n1918# 0.66fF
C138 a_664_n251# g1 0.18fF
C139 vddc4 a_659_n1911# 0.81fF
C140 w_644_n126# c0 0.06fF
C141 p4 a_659_n1911# 0.08fF
C142 g3 a_652_n2046# 0.04fF
C143 vddc3 c3 0.44fF
C144 gndc4 a_641_n2188# 0.55fF
C145 p3 a_634_n1180# 0.15fF
C146 g1 a_681_n251# 0.19fF
C147 a_652_n2046# c0 0.09fF
C148 g4 g1 0.09fF
C149 g4 p1 0.09fF
C150 w_626_n700# p2 0.42fF
C151 GG a_652_n2046# 0.09fF
C152 a_606_n2188# a_641_n2188# 1.03fF
C153 p3 a_652_n2046# 0.09fF
C154 p1 g1 0.56fF
C155 p4 c0 0.10fF
C156 a_678_n2188# w_538_n1918# 1.15fF
C157 a_653_n1431# c3 0.05fF
C158 GG p4 0.09fF
C159 p3 p4 0.09fF
C160 a_561_n1431# a_579_n1432# 0.82fF
C161 vddc1 a_681_n251# 0.02fF
C162 vddc3 a_653_n1431# 0.03fF
C163 vddc2 a_639_n692# 2.46fF
C164 GG a_688_n831# 0.18fF
C165 a_652_n2046# w_538_n1918# 0.07fF
C166 vddc4 a_588_n1911# 1.86fF
C167 vddc4 w_538_n1918# 1.22fF
C168 gndc3 c3 0.21fF
C169 c4 Gnd 0.92fF
C170 a_678_n2188# Gnd 2.61fF
C171 a_641_n2188# Gnd 0.33fF
C172 a_606_n2188# Gnd 0.33fF
C173 a_623_n1911# Gnd 0.00fF
C174 a_570_n2188# Gnd 0.35fF
C175 a_551_n2188# Gnd 0.24fF
C176 gndc4 Gnd 1.03fF
C177 a_588_n1911# Gnd 0.03fF
C178 a_551_n1911# Gnd 0.02fF
C179 vddc4 Gnd 0.34fF
C180 g4 Gnd 2.85fF
C181 p4 Gnd 2.54fF
C182 a_652_n2046# Gnd 3.37fF
C183 c3 Gnd 1.02fF
C184 a_653_n1431# Gnd 2.16fF
C185 a_615_n1432# Gnd 0.30fF
C186 a_634_n1180# Gnd 0.13fF
C187 a_579_n1432# Gnd 0.30fF
C188 a_561_n1431# Gnd 0.19fF
C189 gndc3 Gnd 1.21fF
C190 a_561_n1181# Gnd 0.09fF
C191 vddc3 Gnd 0.46fF
C192 g3 Gnd 2.76fF
C193 p3 Gnd 5.94fF
C194 a_651_n831# Gnd 0.27fF
C195 gndc2 Gnd 1.70fF
C196 c2 Gnd 0.23fF
C197 a_688_n831# Gnd 0.85fF
C198 GG Gnd 8.02fF
C199 p2 Gnd 7.26fF
C200 vddc2 Gnd 0.44fF
C201 a_664_n251# Gnd 0.10fF
C202 gndc1 Gnd 0.64fF
C203 c1 Gnd 0.53fF
C204 a_681_n251# Gnd 1.41fF
C205 a_664_n120# Gnd 0.06fF
C206 vddc1 Gnd 0.24fF
C207 g1 Gnd 9.25fF
C208 p1 Gnd 8.22fF
C209 c0 Gnd 6.96fF
C210 w_538_n1918# Gnd 45.34fF
C211 w_545_n1187# Gnd 34.45fF
C212 w_626_n700# Gnd 19.38fF
C213 w_644_n126# Gnd 10.46fF


.tran 0.1n 40n

.control


run
set curplottitle="Sanjana Sheela - 20231012027- postlayout"
plot v(c0) v(c1)+2 v(c2)+4 (c3)+6 v(c4)+8
plot v(p1) v(g1)+2 v(c0)+4 v(c1)+6
plot v(p2) v(g2)+2 v(c1)+4 v(c2)+6
plot v(p3) v(g3)+2 v(c2)+4 v(c3)+6
plot v(p4) v(g4)+2 v(c3)+4 v(c4)+6

.endc
.end


* postlayout
.include TSMC_180nm.txt
.param LAMBDA=0.09u
.param SUPPLY=1.8
.param width=1.8n
.param width_P=2*width
.param width_N=width
.global gnd vdd

VD1 vdd1 0 1.8V
VD2 vdd11 0 1.8V
VD3 vdd2 0 1.8V
VD4 vdd22 0 1.8V
VD5 vddc1 0 1.8V
VD6 vddc2 0 1.8V
VD7 vdd33 0 1.8V
VD8 vdd3 0 1.8V
VD9 vddc3 0 1.8V
VD10 vdd44 0 1.8V
VD11 vdd4 0 1.8V
VD12 vddc4 0 1.8V
VD13 vdds1 0 1.8V
VD14 vdds2 0 1.8V
VD15 vdds3 0 1.8V
VD16 vdds4 0 1.8V


VG1 gnd1 0 0
VG2 gnd11 0 0
VG3 gnd2 0 0
VG4 gnd22 0 0
VG5 gndc2 0 0
VG6 gndc1 0 0
VG7 gnd3 0 0
VG8 gnd33 0 0
VG9 gndc3 0 0
VG10 gnd4 0 0
VG11 gnd44 0 0
VG12 gndc4 0 0
VG13 gnds1 0 0
VG14 gnds2 0 0
VG15 gnds3 0 0
VG16 gnds4 0 0

VDD vdd gnd 'SUPPLY'

Va1 a1i gnd pulse(0 0 1n 0 0 1n 2n)
Va2 a2i gnd pulse(0 0 1n 0 0 2n 4n)
Va3 a3i gnd pulse(0 0 1n 0 0 4n 8n)
Va4 a4i gnd pulse(0 0 1n 0 0 8n 16n)

Vb4 b4i gnd pulse(1.8 1.8 1n 0 0 16n 32n)
Vb3 b3i gnd pulse(1.8 1.8 1n 0 0 32n 64n)
Vb2 b2i gnd pulse(1.8 1.8 1n 0 0 64n 128n)
Vb1 b1i gnd pulse(1.8 1.8 1n 0 0 128n 256n)

Vcin c0i gnd pulse(0 0 1n 0 0 1n 2n)

Vclk clk gnd pulse(0 1.8 0.2n 0 0 0.5n 1n)

* Va1 b4i gnd pulse(1.8 0 1n 0 0 10n 20n)
* Va2 b3i gnd pulse(1.8 0 1n 0 0 20n 40n)
* Va3 b2i gnd pulse(1.8 0 1n 0 0 40n 80n)
* Va4 b1i gnd pulse(1.8 0 1n 0 0 80n 160n)

* Vb4 a4i gnd pulse(1.8 0 1n 0 0 160n 320n)
* Vb3 a3i gnd pulse(1.8 0 1n 0 0 320n 640n)
* Vb2 a2i gnd pulse(1.8 0 1n 0 0 640n 1280n)
* Vb1 a1i gnd pulse(1.8 0 1n 0 0 1280n 2560n)

* Vcin c0i gnd pulse(1.8 0 1n 0 0 5n 10n)

* Vclk clk gnd pulse(0 1.8 0.2n 0 0 5n 10n)



.option scale=0.09u

M1000 a_1131_n563# s3o vdd w_1124_n466# CMOSP w=40 l=2
+  ad=200 pd=90 as=17870 ps=8038
M1001 a_725_n1062# p4 gnds4 Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=95 ps=48
M1002 gndc2 g1 a_529_n630# Gnd CMOSN w=30 l=2
+  ad=650 pd=300 as=750 ps=330
M1003 vddc4 p1 a_506_n1355# w_493_n1362# CMOSP w=200 l=2
+  ad=3280 pd=1372 as=3000 ps=1230
M1004 vdd a_n184_n277# a_n93_n282# w_n7_n341# CMOSP w=40 l=2
+  ad=0 pd=0 as=395 ps=178
M1005 gnd a_n99_n79# a_n76_n145# Gnd CMOSN w=20 l=2
+  ad=8900 pd=4450 as=200 ps=100
M1006 a_168_n623# b2 vdd22 w_162_n557# CMOSP w=40 l=2
+  ad=400 pd=180 as=600 ps=270
M1007 a_964_n564# a_913_n631# vdd w_849_n466# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1008 a_958_n630# clk a_964_n564# Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=100 ps=50
M1009 a_608_n1088# p3 a_570_n1089# Gnd CMOSN w=80 l=2
+  ad=500 pd=220 as=930 ps=402
M1010 a_799_n1491# clk a_802_n1315# w_798_n1426# CMOSP w=39 l=2
+  ad=195 pd=88 as=395 ps=178
M1011 c0 a_394_47# gnd Gnd CMOSN w=20 l=2
+  ad=195 pd=98 as=0 ps=0
M1012 gnd a_789_n2# a_849_n2# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1013 gnd a_71_n1682# a_201_n1677# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1014 a_561_n1632# p2 a_525_n1632# Gnd CMOSN w=100 l=2
+  ad=1165 pd=496 as=1250 ps=530
M1015 b1 a_93_26# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1016 a_913_n297# clk a_913_n230# Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=100 ps=50
M1017 s3 p3 c2 Vdd CMOSP w=40 l=2
+  ad=400 pd=180 as=400 ps=180
M1018 gndc3 g1 a_534_n1089# Gnd CMOSN w=40 l=2
+  ad=930 pd=422 as=1000 ps=430
M1019 p4 a4 a_172_n1419# Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=190 ps=96
M1020 gnd a_779_n298# a_839_n298# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1021 gnd33 b3 a_175_n1052# Gnd CMOSN w=40 l=2
+  ad=300 pd=140 as=400 ps=180
M1022 a_890_n1423# a_873_n1423# vdd w_735_n1326# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1023 vdd a_394_47# c0 w_492_96# CMOSP w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1024 s4 a_725_n1062# c3 Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=195 ps=98
M1025 gnd a_997_n991# s4o Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1026 gnd a_69_n1734# a_71_n1682# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1027 c4 a_633_n1632# vddc4 w_493_n1362# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1028 gndc4 g1 a_525_n1632# Gnd CMOSN w=50 l=2
+  ad=1240 pd=556 as=0 ps=0
M1029 a_n99_n1099# a_n99_n1116# vdd w_n105_n1259# CMOSP w=41 l=2
+  ad=205 pd=92 as=0 ps=0
M1030 gndc3 g2 a_570_n1089# Gnd CMOSN w=26 l=2
+  ad=0 pd=0 as=0 ps=0
M1031 a_906_n1059# clk a_909_n883# w_905_n994# CMOSP w=39 l=2
+  ad=195 pd=88 as=395 ps=178
M1032 gndc4 g3 a_596_n1632# Gnd CMOSN w=25 l=2
+  ad=0 pd=0 as=1125 ps=480
M1033 vdd c0i a_400_222# w_492_96# CMOSP w=40 l=2
+  ad=0 pd=0 as=395 ps=178
M1034 a_169_n461# b2 vdd2 w_154_n425# CMOSP w=40 l=2
+  ad=200 pd=90 as=200 ps=90
M1035 a_26_n947# clk a_26_n880# Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=100 ps=50
M1036 a_589_n837# g2 a_552_n838# w_500_n844# CMOSP w=160 l=2
+  ad=1870 pd=778 as=2000 ps=830
M1037 a_802_n1315# a_739_n1491# vdd w_735_n1326# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 vdd a_14_139# a_105_134# w_191_75# CMOSP w=40 l=2
+  ad=0 pd=0 as=395 ps=178
M1039 s1 a_673_n77# c0 Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=0 ps=0
M1040 a_n99_n215# clk a_n184_n277# w_n111_n233# CMOSP w=39 l=2
+  ad=395 pd=178 as=195 ps=88
M1041 p2 b2 a2 w_196_n392# CMOSP w=40 l=2
+  ad=600 pd=270 as=400 ps=180
M1042 gnd a_850_n1424# a_873_n1490# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1043 a_873_n1490# clk a_873_n1423# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1044 gnd a_n110_n1558# a_n50_n1558# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1045 a_566_n630# g2 a_548_n492# w_504_n499# CMOSP w=120 l=2
+  ad=600 pd=250 as=1500 ps=630
M1046 a_n96_n1244# b3i vdd w_n105_n1259# CMOSP w=40 l=2
+  ad=395 pd=178 as=0 ps=0
M1047 a_393_69# clk a_330_88# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=200 ps=100
M1048 a_92_48# clk a_29_67# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=200 ps=100
M1049 g1 a_146_n309# vdd1 w_140_n243# CMOSP w=40 l=2
+  ad=200 pd=90 as=600 ps=270
M1050 a_n65_n493# a_n128_n669# vdd w_n132_n504# CMOSP w=40 l=2
+  ad=395 pd=178 as=0 ps=0
M1051 vddc3 p3 a_589_n837# w_500_n844# CMOSP w=54 l=2
+  ad=2470 pd=1038 as=0 ps=0
M1052 s4 p4 c3 Vdd CMOSP w=40 l=2
+  ad=400 pd=180 as=400 ps=180
M1053 a_201_n1677# clk a_69_n1656# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1054 gnd a_n50_n1558# a_n5_n1557# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1055 gnd a_24_n1490# a_41_n1490# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1056 gnd a_799_n1491# a_844_n1490# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1057 a_1_n1491# a_n50_n1558# vdd w_n114_n1393# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1058 a_400_222# clk a_315_160# w_388_204# CMOSP w=39 l=2
+  ad=0 pd=0 as=195 ps=88
M1059 p3 a3 a_169_n890# Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=190 ps=96
M1060 gnd s4o a_1131_n991# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1061 a_633_n1632# p4 a_596_n1632# Gnd CMOSN w=100 l=2
+  ad=600 pd=260 as=0 ps=0
M1062 g2 a_168_n623# vdd22 w_162_n557# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1063 vddc2 p2 a_548_n492# w_504_n499# CMOSP w=60 l=2
+  ad=1700 pd=720 as=0 ps=0
M1064 a_172_n1419# b4 vdd4 w_158_n1387# CMOSP w=40 l=2
+  ad=200 pd=90 as=200 ps=90
M1065 gnd b3i a_n99_n1194# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1066 gnd a_980_n991# a_997_n991# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1067 a_n23_n668# clk a_n17_n602# Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=100 ps=50
M1068 a_517_n630# c0 gndc2 Gnd CMOSN w=60 l=2
+  ad=600 pd=140 as=0 ps=0
M1069 gnd a_739_n1491# a_799_n1491# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1070 a_171_n1581# a4 vdd44 w_165_n1515# CMOSP w=40 l=2
+  ad=400 pd=180 as=600 ps=270
M1071 a_n110_n1487# a4i vdd w_n114_n1393# CMOSP w=40 l=2
+  ad=395 pd=178 as=0 ps=0
M1072 vdd a2i a_n99_n215# w_n7_n341# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1073 gnd s2 a_779_n298# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1074 gnd a_1004_n563# s3o Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1075 vdd a_315_160# a_406_155# w_492_96# CMOSP w=40 l=2
+  ad=0 pd=0 as=395 ps=178
M1076 a_894_n1# clk a_900_65# Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=100 ps=50
M1077 a_146_n309# a1 vdd1 w_140_n243# CMOSP w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1078 a_548_n492# g1 a_517_n491# w_504_n499# CMOSP w=120 l=2
+  ad=0 pd=0 as=1800 ps=510
M1079 a_913_n631# clk a_916_n455# w_912_n566# CMOSP w=39 l=2
+  ad=195 pd=88 as=395 ps=178
M1080 gnd a_913_n631# a_958_n630# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1081 s1 c0 a_673_n77# Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=190 ps=96
M1082 gndc4 g4 a_633_n1632# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1083 a_873_n1423# a_850_n1424# vdd w_735_n1326# CMOSP w=41 l=2
+  ad=205 pd=92 as=0 ps=0
M1084 a_739_n1491# clk a_739_n1420# w_731_n1432# CMOSP w=39 l=2
+  ad=195 pd=88 as=395 ps=178
M1085 a2 a_n105_n390# gnd Gnd CMOSN w=20 l=2
+  ad=195 pd=98 as=0 ps=0
M1086 a_168_n623# a2 vdd22 w_162_n557# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 gnd b4i a_69_n1734# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1088 a_n96_n1192# a_n99_n1194# vdd w_n105_n1259# CMOSP w=40 l=2
+  ad=395 pd=178 as=0 ps=0
M1089 gnd a_6_n601# a_23_n601# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1090 a_171_n1581# b4 vdd44 w_165_n1515# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1091 a_n48_n948# clk a_n45_n772# w_n49_n883# CMOSP w=39 l=2
+  ad=195 pd=88 as=395 ps=178
M1092 gnd s2o a_1064_n230# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1093 b2 a_23_n601# vdd w_n132_n504# CMOSP w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1094 a_566_n630# p2 a_529_n630# Gnd CMOSN w=60 l=2
+  ad=400 pd=180 as=0 ps=0
M1095 gndc2 g2 a_566_n630# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1096 gnd b2i a_n128_n669# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1097 c1 a_529_n251# gndc1 Gnd CMOSN w=20 l=2
+  ad=195 pd=98 as=400 ps=190
M1098 p1 a_147_n147# a1 Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=195 ps=98
M1099 a_n97_n1142# clk a_n96_n1192# w_n5_n1196# CMOSP w=39 l=2
+  ad=195 pd=88 as=0 ps=0
M1100 s2 c1 p2 Vdd CMOSP w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1101 a_69_n1617# a_69_n1639# vdd w_63_n1799# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1102 gnd44 a_171_n1581# g4 Gnd CMOSN w=20 l=2
+  ad=300 pd=140 as=100 ps=50
M1103 a_n59_n78# a_n76_n78# vdd w_n214_19# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1104 a_147_n147# b1 gnd11 Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=95 ps=48
M1105 c4o a_890_n1423# vdd w_735_n1326# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1106 a_900_65# a_849_n2# vdd w_785_163# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1107 a_71_n1682# clk a_72_n1732# w_163_n1736# CMOSP w=39 l=2
+  ad=195 pd=88 as=395 ps=178
M1108 a_41_n1490# a_24_n1490# vdd w_n114_n1393# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1109 a_n147_30# a_n210_n146# vdd w_n214_19# CMOSP w=40 l=2
+  ad=395 pd=178 as=0 ps=0
M1110 a_529_n251# p1 a_512_n251# Gnd CMOSN w=40 l=2
+  ad=300 pd=140 as=400 ps=180
M1111 a_n5_n1557# clk a_1_n1491# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1112 gnd s1 a_789_n2# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1113 a_169_n461# b2 gnd2 Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=95 ps=48
M1114 gnd a_849_n2# a_894_n1# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 a_n17_n602# a_n68_n669# vdd w_n132_n504# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1116 a_169_n890# b3 vdd3 w_155_n858# CMOSP w=40 l=2
+  ad=200 pd=90 as=200 ps=90
M1117 vddc4 p2 a_543_n1355# w_493_n1362# CMOSP w=100 l=2
+  ad=0 pd=0 as=2500 ps=1030
M1118 a_543_n1355# g1 a_506_n1355# w_493_n1362# CMOSP w=200 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 gnd a_n99_n1099# a_n99_n1077# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1120 a_779_n298# clk a_779_n227# w_771_n239# CMOSP w=39 l=2
+  ad=195 pd=88 as=395 ps=178
M1121 a_529_n630# p1 a_517_n630# Gnd CMOSN w=60 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 gndc3 g3 a_608_n1088# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 c3 a_608_n1088# gndc3 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 a_614_n1355# g3 a_578_n1355# w_493_n1362# CMOSP w=200 l=2
+  ad=2250 pd=930 as=2330 ps=962
M1125 vddc4 p3 a_578_n1355# w_493_n1362# CMOSP w=66 l=2
+  ad=0 pd=0 as=0 ps=0
M1126 p4 a_172_n1419# a4 Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=195 ps=98
M1127 s3 a_734_n545# c2 Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=195 ps=98
M1128 a_n128_n669# clk a_n128_n598# w_n136_n610# CMOSP w=39 l=2
+  ad=195 pd=88 as=395 ps=178
M1129 a_n169_n349# a_n184_n351# gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1130 a_734_n545# p3 gnds3 Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=95 ps=48
M1131 a_909_n883# a_846_n1059# vdd w_842_n894# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1132 a_n128_n598# b2i vdd w_n132_n504# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1133 gnd a_853_n631# a_913_n631# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1134 gnd s4 a_846_n1059# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1135 a_315_86# clk a_330_117# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=200 ps=100
M1136 a_1053_66# s1o vdd w_1046_163# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1137 gnd a_930_n230# s2o Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1138 p2 a2 b2 w_196_n392# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1139 c3 a_608_n1088# vddc3 w_500_n844# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 gnd a_n76_n78# a_n59_n78# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1141 a_n184_n351# clk a_n169_n320# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=200 ps=100
M1142 a_516_n838# c0 vddc3 w_500_n844# CMOSP w=160 l=2
+  ad=2400 pd=990 as=0 ps=0
M1143 vddc3 p2 a_552_n838# w_500_n844# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1144 gnd a_1_n1491# a_24_n1557# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1145 p3 b3 a3 w_198_n821# CMOSP w=40 l=2
+  ad=600 pd=270 as=400 ps=180
M1146 s4 c3 p4 Vdd CMOSP w=40 l=2
+  ad=0 pd=0 as=600 ps=270
M1147 a_69_n1656# a_71_n1682# vdd w_63_n1799# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1148 a_330_88# a_315_86# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1149 gnd a_957_n992# a_980_n1058# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1150 a_n50_n1558# clk a_n47_n1382# w_n51_n1493# CMOSP w=39 l=2
+  ad=195 pd=88 as=395 ps=178
M1151 a_14_65# clk a_29_96# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=200 ps=100
M1152 a_658_n289# p2 gnds2 Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=95 ps=48
M1153 a_16_94# a_14_139# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1154 a_673_n77# p1 gnds1 Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=95 ps=48
M1155 gnd a_43_n880# a3 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=195 ps=98
M1156 a_1064_n230# s2o vdd w_1057_n133# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1157 a_n45_n772# a_n108_n948# vdd w_n112_n783# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1158 gnd1 a_146_n309# g1 Gnd CMOSN w=20 l=2
+  ad=300 pd=140 as=100 ps=50
M1159 gnd a_906_n1059# a_951_n1058# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1160 gnd a_n99_n1116# a_32_n1114# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1161 a1 a_n59_n78# vdd w_n214_19# CMOSP w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1162 a_24_n1490# a_1_n1491# vdd w_n114_n1393# CMOSP w=41 l=2
+  ad=205 pd=92 as=0 ps=0
M1163 a_29_67# a_14_65# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1164 a_n105_n390# a_n106_n368# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1165 a_516_n1088# c0 gndc3 Gnd CMOSN w=80 l=2
+  ad=800 pd=340 as=0 ps=0
M1166 a_534_n1089# p1 a_516_n1088# Gnd CMOSN w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 a_633_n1632# g4 a_614_n1355# w_493_n1362# CMOSP w=200 l=2
+  ad=1000 pd=410 as=0 ps=0
M1168 a_846_n1059# clk a_846_n988# w_838_n1000# CMOSP w=39 l=2
+  ad=195 pd=88 as=395 ps=178
M1169 gnd a_41_n1490# a4 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 a_529_n251# g1 a_512_n120# w_492_n126# CMOSP w=80 l=2
+  ad=400 pd=170 as=1200 ps=510
M1171 gnd a_913_n230# a_930_n230# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1172 a_916_n455# a_853_n631# vdd w_849_n466# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1173 gnd33 a_168_n1052# g3 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1174 c4 a_633_n1632# gndc4 Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1175 gnd c4o a_1024_n1423# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1176 s2 a_658_n289# c1 Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=0 ps=0
M1177 gnd s3 a_853_n631# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1178 a_178_n1581# a4 a_171_n1581# Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=200 ps=90
M1179 vdd a_92_48# a_93_26# w_191_75# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1180 a_n184_n277# a2i gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1181 s4o a_997_n991# vdd w_842_n894# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1182 gnd a_n59_n78# a1 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1183 vddc1 p1 a_512_n120# w_492_n126# CMOSP w=80 l=2
+  ad=1000 pd=430 as=0 ps=0
M1184 vddc3 p1 a_516_n838# w_500_n844# CMOSP w=160 l=2
+  ad=0 pd=0 as=0 ps=0
M1185 s1 c0 p1 Vdd CMOSP w=40 l=2
+  ad=400 pd=180 as=600 ps=270
M1186 b4 a_69_n1617# vdd w_63_n1799# CMOSP w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1187 vdd a_n182_n322# a_n184_n351# w_n7_n341# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1188 vdd a_n184_n351# a_n106_n368# w_n7_n341# CMOSP w=41 l=2
+  ad=0 pd=0 as=205 ps=92
M1189 a_517_n491# c0 vddc2 w_504_n499# CMOSP w=120 l=2
+  ad=0 pd=0 as=0 ps=0
M1190 gnd a_987_n563# a_1004_n563# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1191 a_168_n1052# b3 vdd33 w_162_n986# CMOSP w=40 l=2
+  ad=400 pd=180 as=600 ps=270
M1192 vdd a_n105_n390# a2 w_n7_n341# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1193 gnd44 b4 a_178_n1581# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 gnd a4i a_n110_n1558# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1195 a_850_n1424# a_799_n1491# vdd w_735_n1326# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1196 a_890_n231# a_839_n298# vdd w_775_n133# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1197 s2o a_930_n230# vdd w_775_n133# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1198 a_884_n297# clk a_890_n231# Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=100 ps=50
M1199 a_n76_n145# clk a_n76_n78# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1200 gnd a3i a_n108_n948# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1201 gnd a_n99_n1077# b3 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1202 a_1131_n991# s4o vdd w_1124_n894# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1203 a_14_139# b1i gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1204 a_6_n668# clk a_6_n601# Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=100 ps=50
M1205 gnd a_n17_n602# a_6_n668# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1206 a_997_n991# a_980_n991# vdd w_842_n894# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1207 a_24_n1557# clk a_24_n1490# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1208 a_n150_n146# clk a_n147_30# w_n151_n81# CMOSP w=39 l=2
+  ad=195 pd=88 as=0 ps=0
M1209 a3 a_43_n880# vdd w_n112_n783# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1210 a_69_n1639# a_69_n1656# vdd w_63_n1799# CMOSP w=41 l=2
+  ad=205 pd=92 as=0 ps=0
M1211 p4 a4 b4 w_201_n1350# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 a_23_n601# a_6_n601# vdd w_n132_n504# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1213 gndc4 g2 a_561_n1632# Gnd CMOSN w=33 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 a_n210_n75# a1i vdd w_n214_19# CMOSP w=40 l=2
+  ad=395 pd=178 as=0 ps=0
M1215 s3o a_1004_n563# vdd w_849_n466# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1216 gnd s3o a_1131_n563# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1217 a_980_n1058# clk a_980_n991# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1218 gnd a_69_n1639# a_69_n1617# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1219 a_317_115# a_315_160# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1220 s1o a_940_66# vdd w_785_163# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1221 gnd1 b1 a_153_n309# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1222 a_552_n838# g1 a_516_n838# w_500_n844# CMOSP w=160 l=2
+  ad=0 pd=0 as=0 ps=0
M1223 vdd a_14_65# a_92_48# w_191_75# CMOSP w=41 l=2
+  ad=0 pd=0 as=205 ps=92
M1224 a_849_n2# clk a_852_174# w_848_63# CMOSP w=39 l=2
+  ad=195 pd=88 as=395 ps=178
M1225 a_n108_n877# a3i vdd w_n112_n783# CMOSP w=40 l=2
+  ad=395 pd=178 as=0 ps=0
M1226 a_330_117# a_317_115# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 a_6_n601# a_n17_n602# vdd w_n132_n504# CMOSP w=41 l=2
+  ad=205 pd=92 as=0 ps=0
M1228 a_72_n1784# b4i vdd w_63_n1799# CMOSP w=40 l=2
+  ad=395 pd=178 as=0 ps=0
M1229 a4 a_41_n1490# vdd w_n114_n1393# CMOSP w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1230 a_930_n230# a_913_n230# vdd w_775_n133# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1231 p2 a_169_n461# a2 Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=0 ps=0
M1232 g3 a_168_n1052# vdd33 w_162_n986# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1233 a_n110_n1558# clk a_n110_n1487# w_n118_n1499# CMOSP w=39 l=2
+  ad=195 pd=88 as=0 ps=0
M1234 a_n182_n322# a_n184_n277# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1235 gnd22 b2 a_175_n623# Gnd CMOSN w=40 l=2
+  ad=300 pd=140 as=400 ps=180
M1236 a_512_n251# c0 gndc1 Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1237 a_n99_n79# a_n150_n146# vdd w_n214_19# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1238 gnd a_n128_n669# a_n68_n669# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1239 a_n108_n948# clk a_n108_n877# w_n116_n889# CMOSP w=39 l=2
+  ad=195 pd=88 as=0 ps=0
M1240 gnd a_873_n1423# a_890_n1423# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1241 p1 a1 b1 w_176_n77# CMOSP w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1242 a_n93_n282# clk a_n182_n322# w_n105_n300# CMOSP w=39 l=2
+  ad=0 pd=0 as=195 ps=88
M1243 a_608_n1088# g3 a_589_n837# w_500_n844# CMOSP w=160 l=2
+  ad=800 pd=330 as=0 ps=0
M1244 gnd a_69_n1656# a_200_n1654# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1245 s3 c2 p3 Vdd CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1246 p3 a3 b3 w_198_n821# CMOSP w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1247 c1 a_529_n251# vddc1 w_492_n126# CMOSP w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1248 gnd a_n68_n669# a_n23_n668# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1249 a_951_n1058# clk a_957_n992# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1250 a_172_n1419# b4 gnd4 Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=95 ps=48
M1251 a_32_n1114# clk a_n99_n1099# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1252 vddc2 p1 a_517_n491# w_504_n499# CMOSP w=120 l=2
+  ad=0 pd=0 as=0 ps=0
M1253 a_779_n227# s2 vdd w_775_n133# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1254 a_105_134# clk a_16_94# w_93_116# CMOSP w=39 l=2
+  ad=0 pd=0 as=195 ps=88
M1255 gnd a_940_66# s1o Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1256 a_839_n298# clk a_842_n122# w_838_n233# CMOSP w=39 l=2
+  ad=195 pd=88 as=395 ps=178
M1257 gnd22 a_168_n623# g2 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1258 a_987_n630# clk a_987_n563# Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=100 ps=50
M1259 a_168_n1052# a3 vdd33 w_162_n986# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1260 a_980_n991# a_957_n992# vdd w_842_n894# CMOSP w=41 l=2
+  ad=205 pd=92 as=0 ps=0
M1261 gnd a_846_n1059# a_906_n1059# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1262 a_506_n1632# c0 gndc4 Gnd CMOSN w=100 l=2
+  ad=1000 pd=420 as=0 ps=0
M1263 a_940_66# a_923_66# vdd w_785_163# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1264 vdd a_93_26# b1 w_191_75# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1265 a_570_n1089# p2 a_534_n1089# Gnd CMOSN w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1266 a_844_n1490# clk a_850_n1424# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1267 a_n99_n1077# a_n99_n1099# vdd w_n105_n1259# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1268 vdd a_16_94# a_14_65# w_191_75# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1269 s2 c1 a_658_n289# Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=0 ps=0
M1270 gnd a_26_n880# a_43_n880# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1271 a_789_n2# clk a_789_69# w_781_57# CMOSP w=39 l=2
+  ad=195 pd=88 as=395 ps=178
M1272 gnd a1i a_n210_n146# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1273 vdd a_n106_n368# a_n105_n390# w_n7_n341# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1274 gnd a_964_n564# a_987_n630# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1275 a_525_n1632# p1 a_506_n1632# Gnd CMOSN w=100 l=2
+  ad=0 pd=0 as=0 ps=0
M1276 a_72_n1732# a_69_n1734# vdd w_63_n1799# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1277 a_n76_n78# a_n99_n79# vdd w_n214_19# CMOSP w=41 l=2
+  ad=205 pd=92 as=0 ps=0
M1278 a_725_n1062# p4 vdds4 Vdd CMOSP w=40 l=2
+  ad=200 pd=90 as=200 ps=90
M1279 a_153_n309# a1 a_146_n309# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1280 a_n47_n1382# a_n110_n1558# vdd w_n114_n1393# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1281 a_406_155# clk a_317_115# w_394_137# CMOSP w=39 l=2
+  ad=0 pd=0 as=195 ps=88
M1282 c2 a_566_n630# gndc2 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1283 a_169_n890# b3 gnd3 Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=95 ps=48
M1284 s4 c3 a_725_n1062# Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=0 ps=0
M1285 a_315_160# c0i gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1286 p1 b1 a1 w_176_n77# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1287 gnd a_890_n231# a_913_n297# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1288 a_987_n563# a_964_n564# vdd w_849_n466# CMOSP w=41 l=2
+  ad=205 pd=92 as=0 ps=0
M1289 a_739_n1420# c4 vdd w_735_n1326# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1290 a_394_47# a_393_69# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1291 a_147_n147# b1 vdd11 w_134_n112# CMOSP w=40 l=2
+  ad=200 pd=90 as=200 ps=90
M1292 a_853_n631# clk a_853_n560# w_845_n572# CMOSP w=39 l=2
+  ad=195 pd=88 as=395 ps=178
M1293 gnd a_n97_n1142# a_33_n1137# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1294 a_93_26# a_92_48# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1295 gndc1 g1 a_529_n251# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1296 a_175_n623# a2 a_168_n623# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1297 gnd c4 a_739_n1491# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1298 a_29_96# a_16_94# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1299 a_512_n120# c0 vddc1 w_492_n126# CMOSP w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1300 a_846_n988# s4 vdd w_842_n894# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1301 a_578_n1355# g2 a_543_n1355# w_493_n1362# CMOSP w=200 l=2
+  ad=0 pd=0 as=0 ps=0
M1302 gnd a_69_n1617# b4 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1303 vdd a_393_69# a_394_47# w_492_96# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1304 a_3_n881# a_n48_n948# vdd w_n112_n783# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1305 a_n3_n947# clk a_3_n881# Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=100 ps=50
M1306 a_69_n1734# clk a_72_n1784# w_169_n1803# CMOSP w=39 l=2
+  ad=195 pd=88 as=0 ps=0
M1307 a_n99_n1194# clk a_n96_n1244# w_1_n1263# CMOSP w=39 l=2
+  ad=195 pd=88 as=0 ps=0
M1308 a_923_66# a_900_65# vdd w_785_163# CMOSP w=41 l=2
+  ad=205 pd=92 as=0 ps=0
M1309 gnd a_900_65# a_923_n1# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1310 gnd a_n150_n146# a_n105_n145# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1311 p4 b4 a4 w_201_n1350# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1312 vdd a_317_115# a_315_86# w_492_96# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1313 gnd a_923_66# a_940_66# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1314 c2 a_566_n630# vddc2 w_504_n499# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1315 a_n99_n1116# a_n97_n1142# vdd w_n105_n1259# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1316 p3 a_169_n890# a3 Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=0 ps=0
M1317 gnd a_890_n1423# c4o Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1318 p1 a1 a_147_n147# Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=0 ps=0
M1319 a_734_n545# p3 vdds3 Vdd CMOSP w=40 l=2
+  ad=200 pd=90 as=200 ps=90
M1320 a_1024_n1423# c4o vdd w_1017_n1326# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1321 a_n105_n145# clk a_n99_n79# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1322 gnd a_n210_n146# a_n150_n146# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1323 a_99_201# clk a_14_139# w_87_183# CMOSP w=39 l=2
+  ad=395 pd=178 as=195 ps=88
M1324 gnd a_23_n601# b2 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1325 a_596_n1632# p3 a_561_n1632# Gnd CMOSN w=100 l=2
+  ad=0 pd=0 as=0 ps=0
M1326 gnd a_839_n298# a_884_n297# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1327 p2 a2 a_169_n461# Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=0 ps=0
M1328 gnd a_3_n881# a_26_n947# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1329 a_200_n1654# clk a_69_n1639# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1330 a_33_n1137# clk a_n99_n1116# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1331 a_923_n1# clk a_923_66# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1332 a_n106_n368# clk a_n169_n349# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1333 a_n210_n146# clk a_n210_n75# w_n218_n87# CMOSP w=39 l=2
+  ad=195 pd=88 as=0 ps=0
M1334 a_913_n230# a_890_n231# vdd w_775_n133# CMOSP w=41 l=2
+  ad=205 pd=92 as=0 ps=0
M1335 a_43_n880# a_26_n880# vdd w_n112_n783# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1336 gnd s1o a_1053_66# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1337 a_957_n992# a_906_n1059# vdd w_842_n894# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1338 a_658_n289# p2 vdds2 Vdd CMOSP w=40 l=2
+  ad=200 pd=90 as=200 ps=90
M1339 a_n68_n669# clk a_n65_n493# w_n69_n604# CMOSP w=39 l=2
+  ad=195 pd=88 as=0 ps=0
M1340 a_1004_n563# a_987_n563# vdd w_849_n466# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1341 a_789_69# s1 vdd w_785_163# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1342 a_852_174# a_789_n2# vdd w_785_163# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1343 a_853_n560# s3 vdd w_849_n466# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1344 vdd b1i a_99_201# w_191_75# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1345 a_673_n77# p1 vdds1 Vdd CMOSP w=40 l=2
+  ad=200 pd=90 as=200 ps=90
M1346 s3 c2 a_734_n545# Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=0 ps=0
M1347 a_26_n880# a_3_n881# vdd w_n112_n783# CMOSP w=41 l=2
+  ad=205 pd=92 as=0 ps=0
M1348 b3 a_n99_n1077# vdd w_n105_n1259# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1349 gnd a_n99_n1194# a_n97_n1142# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1350 gnd a_n108_n948# a_n48_n948# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1351 a_506_n1355# c0 vddc4 w_493_n1362# CMOSP w=200 l=2
+  ad=0 pd=0 as=0 ps=0
M1352 vdd a_315_86# a_393_69# w_492_96# CMOSP w=41 l=2
+  ad=0 pd=0 as=205 ps=92
M1353 a_n169_n320# a_n182_n322# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1354 vddc4 p4 a_614_n1355# w_493_n1362# CMOSP w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1355 g4 a_171_n1581# vdd44 w_165_n1515# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1356 s1 p1 c0 Vdd CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1357 a_842_n122# a_779_n298# vdd w_775_n133# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1358 gnd a_n48_n948# a_n3_n947# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1359 a_146_n309# b1 vdd1 w_140_n243# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1360 s2 p2 c1 Vdd CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1361 a_175_n1052# a3 a_168_n1052# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
C0 a_923_66# w_785_163# 0.17fF
C1 a_16_94# w_93_116# 0.08fF
C2 a_894_n1# clk 0.05fF
C3 a_n17_n602# a_6_n601# 0.05fF
C4 a_14_65# w_191_75# 0.17fF
C5 a1 a_147_n147# 0.05fF
C6 a_1_n1491# a_24_n1490# 0.05fF
C7 g2 p4 0.19fF
C8 a_n108_n948# a_n108_n877# 0.40fF
C9 a_n99_n1116# a_n97_n1142# 0.05fF
C10 a_873_n1490# gnd 0.21fF
C11 b1i a_99_201# 0.05fF
C12 a_789_n2# a_789_69# 0.40fF
C13 a_930_n230# gnd 0.21fF
C14 p1 vdds1 0.03fF
C15 c0 a_673_n77# 0.05fF
C16 w_63_n1799# a_72_n1784# 0.08fF
C17 a_852_174# a_849_n2# 0.40fF
C18 w_775_n133# a_779_n227# 0.08fF
C19 b1i gnd 0.12fF
C20 g2 vdd22 0.44fF
C21 vddc2 a_548_n492# 1.08fF
C22 b3i gnd 0.12fF
C23 a1 a_146_n309# 0.12fF
C24 w_154_n425# b2 0.06fF
C25 a_n99_n79# vdd 0.41fF
C26 w_493_n1362# g1 0.08fF
C27 a_6_n668# gnd 0.21fF
C28 w_1057_n133# s2o 0.09fF
C29 p1 g4 0.09fF
C30 g2 p3 0.41fF
C31 a_93_26# vdd 0.44fF
C32 a_1053_66# gnd 0.23fF
C33 s1o a_1053_66# 0.13fF
C34 c2 p3 0.23fF
C35 a_566_n630# gndc2 0.26fF
C36 w_n7_n341# vdd 0.70fF
C37 a4i a_n110_n1487# 0.05fF
C38 a1i gnd 0.12fF
C39 p2 vdds2 0.03fF
C40 a_850_n1424# a_844_n1490# 0.21fF
C41 a_16_94# a_14_65# 0.05fF
C42 a_853_n631# a_916_n455# 0.05fF
C43 a_41_n1490# vdd 0.44fF
C44 w_849_n466# vdd 0.70fF
C45 w_n114_n1393# a_41_n1490# 0.17fF
C46 a_69_n1639# a_69_n1656# 0.05fF
C47 gnd a_201_n1677# 0.24fF
C48 a_916_n455# a_913_n631# 0.40fF
C49 clk m2_n16_n623# 0.03fF
C50 a_890_n1423# c4o 0.13fF
C51 c0 w_492_96# 0.08fF
C52 w_n112_n783# a3i 0.09fF
C53 b2 vdd 0.44fF
C54 b2 vdd2 0.03fF
C55 w_n214_19# a_n210_n75# 0.08fF
C56 a_n45_n772# a_n48_n948# 0.40fF
C57 gndc4 a_525_n1632# 1.01fF
C58 vddc4 a_543_n1355# 1.86fF
C59 a_n48_n948# a_n3_n947# 0.08fF
C60 a_3_n881# vdd 0.41fF
C61 a_802_n1315# a_799_n1491# 0.40fF
C62 w_n218_n87# clk 0.10fF
C63 b3 a_169_n890# 0.05fF
C64 p3 a_589_n837# 0.15fF
C65 a_315_86# clk 0.02fF
C66 g2 g3 0.29fF
C67 gndc3 a_570_n1089# 0.42fF
C68 w_n214_19# a1 0.08fF
C69 a_1_n1491# a_24_n1557# 0.08fF
C70 g4 a_633_n1632# 0.13fF
C71 a_93_26# gnd 0.21fF
C72 a3i gnd 0.12fF
C73 a_201_n1677# a_71_n1682# 0.08fF
C74 b4 vdd4 0.03fF
C75 a4 a_41_n1490# 0.13fF
C76 w_504_n499# g2 0.07fF
C77 a_14_65# a_92_48# 0.05fF
C78 a_n147_30# a_n150_n146# 0.40fF
C79 a_913_n631# a_958_n630# 0.08fF
C80 c3 a_725_n1062# 0.05fF
C81 a_41_n1490# gnd 0.21fF
C82 a_529_n251# gndc1 0.24fF
C83 w_n112_n783# a_3_n881# 0.17fF
C84 vdd w_191_75# 0.70fF
C85 a3 vdd33 0.02fF
C86 w_504_n499# c2 0.08fF
C87 w_493_n1362# p2 0.66fF
C88 a_799_n1491# clk 0.07fF
C89 w_196_n392# p2 1.63fF
C90 a_779_n298# a_842_n122# 0.05fF
C91 w_165_n1515# vdd44 0.39fF
C92 a_n97_n1142# gnd 0.23fF
C93 a_n96_n1244# vdd 0.44fF
C94 clk m2_4_n902# 0.03fF
C95 a_71_n1682# clk 0.07fF
C96 a_849_n2# a_894_n1# 0.08fF
C97 a_69_n1734# a_72_n1784# 0.40fF
C98 g1 g2 0.42fF
C99 w_735_n1326# c4o 0.08fF
C100 b2 gnd 0.23fF
C101 w_176_n77# b1 0.36fF
C102 a_890_n231# vdd 0.41fF
C103 clk m2_74_90# 0.03fF
C104 s4o a_1131_n991# 0.13fF
C105 a_525_n1632# a_561_n1632# 1.03fF
C106 w_905_n994# clk 0.10fF
C107 a_6_n601# vdd 0.78fF
C108 a_n128_n669# a_n65_n493# 0.05fF
C109 gnd1 b2 0.21fF
C110 a_739_n1420# vdd 0.44fF
C111 c1 a_658_n289# 0.05fF
C112 s2 p2 0.52fF
C113 w_492_n126# c1 0.10fF
C114 a_906_n1059# gnd 0.23fF
C115 p3 a3 0.98fF
C116 a_146_n309# a_153_n309# 0.47fF
C117 a_n128_n669# gnd 0.24fF
C118 w_63_n1799# a_69_n1639# 0.17fF
C119 a_589_n837# a_608_n1088# 1.82fF
C120 w_771_n239# clk 0.10fF
C121 a_29_67# a_92_48# 0.23fF
C122 clk m2_924_46# 0.03fF
C123 p2 a_169_n461# 0.20fF
C124 w_n69_n604# a_n65_n493# 0.07fF
C125 w_n51_n1493# clk 0.10fF
C126 w_842_n894# a_909_n883# 0.08fF
C127 a_171_n1581# vdd44 1.15fF
C128 a_n182_n322# gnd 0.23fF
C129 a_99_201# w_191_75# 0.08fF
C130 s1 w_785_163# 0.09fF
C131 a_844_n1490# gnd 0.24fF
C132 a_842_n122# a_839_n298# 0.40fF
C133 a_849_n2# w_785_163# 0.09fF
C134 c4 a_739_n1420# 0.05fF
C135 p4 a_725_n1062# 0.05fF
C136 a_315_160# a_400_222# 0.40fF
C137 w_162_n986# a3 0.06fF
C138 a_n68_n669# a_n17_n602# 0.05fF
C139 p4 b4 0.52fF
C140 w_1124_n894# s4o 0.09fF
C141 a_n68_n669# a_n23_n668# 0.08fF
C142 a_393_69# w_492_96# 0.17fF
C143 g1 a_529_n630# 0.08fF
C144 a4 vdd44 0.02fF
C145 vdd a_72_n1784# 0.44fF
C146 w_163_n1736# a_71_n1682# 0.08fF
C147 s1 gnd 0.12fF
C148 w_63_n1799# a_72_n1732# 0.08fF
C149 a_997_n991# a_980_n1058# 0.16fF
C150 a_315_160# a_406_155# 0.05fF
C151 p1 vddc1 0.02fF
C152 a_839_n298# a_884_n297# 0.08fF
C153 w_n7_n341# a_n105_n390# 0.17fF
C154 w_905_n994# a_906_n1059# 0.08fF
C155 a_799_n1491# a_844_n1490# 0.08fF
C156 a_849_n2# gnd 0.23fF
C157 w_775_n133# a_930_n230# 0.17fF
C158 a_14_139# a_105_134# 0.05fF
C159 a_178_n1581# gnd44 0.71fF
C160 w_493_n1362# vddc4 1.22fF
C161 p2 g2 1.70fF
C162 a_69_n1639# a_200_n1654# 0.23fF
C163 a_92_48# vdd 0.78fF
C164 a_317_115# a_406_155# 0.40fF
C165 a_16_94# gnd 0.23fF
C166 w_140_n243# a_146_n309# 0.19fF
C167 a_853_n631# gnd 0.24fF
C168 w_n7_n341# a2i 0.09fF
C169 c2 s3 0.98fF
C170 a_957_n992# clk 0.02fF
C171 clk m2_n122_n349# 0.03fF
C172 a_913_n631# gnd 0.23fF
C173 a_330_88# gnd 0.21fF
C174 w_169_n1803# clk 0.10fF
C175 a_n5_n1557# clk 0.05fF
C176 p3 vdds3 0.03fF
C177 s3 a_853_n560# 0.05fF
C178 clk w_394_137# 0.10fF
C179 a_n106_n368# vdd 0.78fF
C180 a_913_n297# gnd 0.21fF
C181 vddc4 a_614_n1355# 0.81fF
C182 a1 vdd1 0.02fF
C183 a_1_n1491# vdd 0.41fF
C184 w_845_n572# clk 0.10fF
C185 w_n214_19# a_n210_n146# 0.09fF
C186 w_n114_n1393# a_1_n1491# 0.17fF
C187 w_154_n425# a_169_n461# 0.06fF
C188 a_29_96# a_14_65# 0.21fF
C189 a_315_86# a_330_88# 0.08fF
C190 vddc1 a_529_n251# 0.02fF
C191 gndc4 a_506_n1632# 1.26fF
C192 vddc4 a_506_n1355# 5.55fF
C193 a_980_n1058# gnd 0.21fF
C194 b1 vdd 0.44fF
C195 a_873_n1490# clk 0.05fF
C196 a_846_n1059# a_909_n883# 0.05fF
C197 a_394_47# w_492_96# 0.17fF
C198 a_n150_n146# gnd 0.23fF
C199 a_516_n1088# a_534_n1089# 0.82fF
C200 w_n151_n81# a_n147_30# 0.07fF
C201 g2 a_570_n1089# 0.08fF
C202 a_n45_n772# vdd 0.44fF
C203 a_6_n668# clk 0.05fF
C204 w_493_n1362# c4 0.54fF
C205 c0 p4 0.21fF
C206 w_781_57# clk 0.10fF
C207 a_26_n880# a_26_n947# 0.23fF
C208 a_n169_n320# a_n184_n351# 0.21fF
C209 a_846_n988# vdd 0.44fF
C210 a_n110_n1558# a_n50_n1558# 0.08fF
C211 vdd a_1024_n1423# 0.44fF
C212 s1 p1 0.52fF
C213 w_838_n233# a_839_n298# 0.08fF
C214 w_n49_n883# clk 0.10fF
C215 p3 a_578_n1355# 0.08fF
C216 w_n214_19# a_n76_n78# 0.17fF
C217 a3 a_168_n1052# 0.12fF
C218 vdd2 a_169_n461# 0.45fF
C219 w_162_n557# a2 0.06fF
C220 a_987_n630# gnd 0.21fF
C221 a_596_n1632# a_633_n1632# 1.03fF
C222 w_176_n77# a1 0.13fF
C223 clk m2_988_n583# 0.03fF
C224 a_n99_n215# vdd 0.44fF
C225 w_504_n499# vddc2 0.75fF
C226 a_201_n1677# clk 0.05fF
C227 w_n132_n504# a_23_n601# 0.17fF
C228 c0 p3 0.39fF
C229 s3o a_1131_n563# 0.13fF
C230 c3 p4 0.21fF
C231 a_906_n1059# a_957_n992# 0.05fF
C232 g1 a_512_n251# 0.18fF
C233 w_n112_n783# a_n45_n772# 0.08fF
C234 w_798_n1426# a_799_n1491# 0.08fF
C235 w_735_n1326# a_890_n1423# 0.17fF
C236 w_492_n126# c0 0.06fF
C237 s4o vdd 0.44fF
C238 w_504_n499# a_548_n492# 0.42fF
C239 w_n7_n341# a_n93_n282# 0.08fF
C240 s2 a_779_n227# 0.05fF
C241 w_838_n1000# clk 0.10fF
C242 a_n128_n669# a_n128_n598# 0.40fF
C243 b1 gnd 0.23fF
C244 a_72_n1732# a_69_n1734# 0.05fF
C245 w_849_n466# a_987_n563# 0.17fF
C246 a_842_n122# vdd 0.44fF
C247 a2 vdd22 0.02fF
C248 a_923_n1# gnd 0.21fF
C249 g4 vdd44 0.44fF
C250 a_997_n991# s4o 0.13fF
C251 w_198_n821# a3 0.13fF
C252 b3 a_n99_n1077# 0.13fF
C253 s2 gnd 0.12fF
C254 a_n99_n1077# vdd 0.44fF
C255 a_n99_n79# clk 0.02fF
C256 w_n118_n1499# clk 0.10fF
C257 a_789_69# vdd 0.44fF
C258 c1 p2 0.53fF
C259 w_492_n126# a_512_n120# 0.35fF
C260 w_63_n1799# b4 0.08fF
C261 w_n114_n1393# a4i 0.09fF
C262 a_n3_n947# gnd 0.24fF
C263 a_1024_n1423# gnd 0.23fF
C264 vdd a_69_n1639# 0.78fF
C265 clk m2_n75_n98# 0.03fF
C266 w_n105_n1259# a_n99_n1116# 0.17fF
C267 a_853_n560# vdd 0.44fF
C268 w_155_n858# vdd3 0.08fF
C269 a_n99_n1194# gnd 0.24fF
C270 g1 a_534_n1089# 0.08fF
C271 w_842_n894# vdd 0.70fF
C272 a_394_47# c0 0.13fF
C273 c0 g3 0.29fF
C274 w_158_n1387# b4 0.09fF
C275 a_400_222# w_492_96# 0.08fF
C276 a_99_201# w_87_183# 0.07fF
C277 b1i w_191_75# 0.09fF
C278 a_32_n1114# a_n99_n1116# 0.08fF
C279 a_n97_n1142# clk 0.07fF
C280 s4o gnd 0.23fF
C281 w_1124_n466# a_1131_n563# 0.08fF
C282 w_162_n557# vdd22 0.39fF
C283 a_789_69# w_785_163# 0.08fF
C284 a_n96_n1244# b3i 0.05fF
C285 a_n182_n322# a_n93_n282# 0.40fF
C286 w_493_n1362# p1 0.08fF
C287 w_n5_n1196# clk 0.10fF
C288 w_504_n499# c0 0.08fF
C289 w_845_n572# a_853_n631# 0.08fF
C290 a_n65_n493# a_n68_n669# 0.40fF
C291 a_406_155# w_492_96# 0.08fF
C292 a_n76_n78# a_n76_n145# 0.23fF
C293 w_842_n894# a_997_n991# 0.17fF
C294 a_n210_n75# vdd 0.44fF
C295 a_739_n1491# gnd 0.24fF
C296 s3o vdd 0.44fF
C297 w_912_n566# a_916_n455# 0.07fF
C298 p1 b1 0.52fF
C299 a_3_n881# clk 0.02fF
C300 vdd a_72_n1732# 0.44fF
C301 a_957_n992# a_980_n1058# 0.08fF
C302 a_315_160# gnd 0.24fF
C303 a_n68_n669# gnd 0.23fF
C304 gndc4 c4 0.24fF
C305 a_608_n1088# c3 0.05fF
C306 c0 g1 0.56fF
C307 a_6_n601# a_6_n668# 0.23fF
C308 a_906_n1059# clk 0.07fF
C309 clk m2_n124_n326# 0.03fF
C310 p3 p4 0.19fF
C311 a_n99_n1077# gnd 0.21fF
C312 w_163_n1736# clk 0.10fF
C313 a_873_n1423# a_890_n1423# 0.18fF
C314 p1 a_506_n1355# 0.08fF
C315 w_n105_n1259# b3 0.08fF
C316 a_n128_n669# clk 0.05fF
C317 w_775_n133# a_890_n231# 0.17fF
C318 a4i gnd 0.12fF
C319 w_n105_n1259# vdd 0.70fF
C320 g2 a_566_n630# 0.18fF
C321 w_140_n243# g1 0.06fF
C322 a_552_n838# a_589_n837# 1.65fF
C323 w_n114_n1393# a_n50_n1558# 0.09fF
C324 a_n106_n368# a_n105_n390# 0.18fF
C325 w_848_63# a_852_174# 0.07fF
C326 a1 vdd 0.44fF
C327 a_n108_n948# a_n48_n948# 0.08fF
C328 a_930_n230# a_913_n297# 0.16fF
C329 a_317_115# gnd 0.23fF
C330 w_162_n986# vdd33 0.39fF
C331 a_566_n630# c2 0.08fF
C332 a_n182_n322# clk 0.07fF
C333 w_500_n844# g2 0.07fF
C334 a_951_n1058# gnd 0.24fF
C335 p2 a_548_n492# 0.08fF
C336 w_n5_n1196# a_n97_n1142# 0.08fF
C337 w_493_n1362# g4 0.07fF
C338 a_844_n1490# clk 0.05fF
C339 a_317_115# a_315_86# 0.05fF
C340 a_29_96# gnd 0.24fF
C341 a_69_n1617# a_69_n1639# 0.18fF
C342 w_169_n1803# a_72_n1784# 0.07fF
C343 a_739_n1491# a_799_n1491# 0.08fF
C344 c2 a_734_n545# 0.05fF
C345 a_884_n297# gnd 0.24fF
C346 w_n69_n604# clk 0.10fF
C347 a_673_n77# gnds1 0.23fF
C348 w_n132_n504# b2i 0.09fF
C349 a_n108_n877# vdd 0.44fF
C350 w_140_n243# vdd1 0.39fF
C351 w_n7_n341# a_n182_n322# 0.09fF
C352 g1 a_146_n309# 0.17fF
C353 s4 a_846_n988# 0.05fF
C354 a_890_n231# clk 0.02fF
C355 a_93_26# w_191_75# 0.17fF
C356 w_493_n1362# a_633_n1632# 1.15fF
C357 a_n110_n1558# a_n47_n1382# 0.05fF
C358 g3 vdd33 0.44fF
C359 s3o gnd 0.23fF
C360 w_n116_n889# clk 0.10fF
C361 w_1124_n466# vdd 0.11fF
C362 w_158_n1387# vdd4 0.08fF
C363 a_1_n1491# a_n5_n1557# 0.21fF
C364 w_n218_n87# a_n210_n75# 0.07fF
C365 a_849_n2# clk 0.07fF
C366 a_614_n1355# a_633_n1632# 2.06fF
C367 a_n96_n1192# vdd 0.44fF
C368 g3 p4 0.19fF
C369 clk m2_965_n585# 0.03fF
C370 a3 b3 0.49fF
C371 a_n210_n146# a_n147_30# 0.05fF
C372 a3 vdd 0.44fF
C373 a_853_n631# clk 0.05fF
C374 a_16_94# clk 0.07fF
C375 c4o vdd 0.44fF
C376 a_168_n623# a_175_n623# 0.47fF
C377 w_798_n1426# a_802_n1315# 0.07fF
C378 a_n50_n1558# gnd 0.23fF
C379 a_n169_n349# gnd 0.21fF
C380 w_735_n1326# a_873_n1423# 0.17fF
C381 w_n112_n783# a_n108_n877# 0.08fF
C382 a1 gnd 0.23fF
C383 a_330_88# clk 0.05fF
C384 a_913_n631# clk 0.07fF
C385 w_n105_n300# a_n93_n282# 0.07fF
C386 a_566_n630# a_529_n630# 0.62fF
C387 p1 g2 0.42fF
C388 w_500_n844# a_589_n837# 0.54fF
C389 a_146_n309# vdd1 1.15fF
C390 a2i a_n99_n215# 0.05fF
C391 a_913_n297# clk 0.05fF
C392 a_32_n1114# gnd 0.21fF
C393 a_516_n838# a_552_n838# 1.65fF
C394 a_n105_n145# gnd 0.24fF
C395 w_n132_n504# a_n17_n602# 0.17fF
C396 p3 g3 0.29fF
C397 c0 p2 0.49fF
C398 a_980_n1058# clk 0.05fF
C399 clk m2_238_n1683# 0.03fF
C400 a_980_n991# vdd 0.78fF
C401 a_393_69# a_394_47# 0.18fF
C402 a_987_n563# a_987_n630# 0.23fF
C403 w_n112_n783# a3 0.08fF
C404 g1 p4 0.19fF
C405 a_534_n1089# a_570_n1089# 0.82fF
C406 vdd w_492_96# 0.70fF
C407 w_849_n466# a_853_n631# 0.09fF
C408 w_n136_n610# a_n128_n598# 0.07fF
C409 a_71_n1682# a_72_n1732# 0.40fF
C410 a_n150_n146# clk 0.07fF
C411 w_798_n1426# clk 0.10fF
C412 w_849_n466# a_913_n631# 0.09fF
C413 a_168_n1052# vdd33 1.15fF
C414 b2 a_168_n623# 0.42fF
C415 a_846_n1059# gnd 0.24fF
C416 w_165_n1515# b4 0.06fF
C417 a_n150_n146# a_n99_n79# 0.05fF
C418 a_923_66# a_923_n1# 0.23fF
C419 a_980_n991# a_997_n991# 0.18fF
C420 w_162_n986# g3 0.06fF
C421 w_134_n112# vdd11 0.08fF
C422 s2o vdd 0.44fF
C423 w_n105_n300# clk 0.10fF
C424 g2 g4 0.09fF
C425 g1 p3 0.38fF
C426 p2 a2 0.99fF
C427 clk m2_n98_n100# 0.03fF
C428 w_842_n894# s4 0.09fF
C429 w_492_n126# g1 0.06fF
C430 b4 vdd 0.44fF
C431 a_169_n461# gnd2 0.22fF
C432 a_n184_n277# gnd 0.24fF
C433 a3 gnd 0.23fF
C434 a_987_n630# clk 0.05fF
C435 a_n99_n1099# a_n99_n1116# 0.05fF
C436 a_940_66# vdd 0.44fF
C437 c4o gnd 0.23fF
C438 w_1017_n1326# vdd 0.11fF
C439 w_n49_n883# a_n45_n772# 0.07fF
C440 w_775_n133# s2 0.09fF
C441 a_n59_n78# a1 0.13fF
C442 a_1_n1491# clk 0.02fF
C443 w_155_n858# b3 0.09fF
C444 c0i w_492_96# 0.09fF
C445 a_92_48# a_93_26# 0.18fF
C446 w_1057_n133# vdd 0.11fF
C447 a1 p1 0.98fF
C448 a_400_222# w_388_204# 0.07fF
C449 g1 a_525_n1632# 0.09fF
C450 a_1004_n563# vdd 0.44fF
C451 w_500_n844# a_516_n838# 0.55fF
C452 w_n51_n1493# a_n50_n1558# 0.08fF
C453 b4 a_171_n1581# 0.42fF
C454 g3 a_608_n1088# 0.17fF
C455 a_957_n992# a_951_n1058# 0.21fF
C456 w_63_n1799# a_69_n1656# 0.17fF
C457 gndc4 a_633_n1632# 0.33fF
C458 a_940_66# w_785_163# 0.17fF
C459 clk m2_914_n250# 0.03fF
C460 a_105_134# w_93_116# 0.07fF
C461 a_16_94# w_191_75# 0.09fF
C462 a_923_n1# clk 0.05fF
C463 a_317_115# w_394_137# 0.08fF
C464 w_n7_n341# a_n106_n368# 0.17fF
C465 s2o a_1064_n230# 0.13fF
C466 w_842_n894# a_957_n992# 0.17fF
C467 w_838_n1000# a_846_n988# 0.07fF
C468 a_n47_n1382# vdd 0.44fF
C469 vddc4 a_578_n1355# 1.13fF
C470 a_n184_n351# vdd 0.41fF
C471 a_315_86# w_492_96# 0.17fF
C472 w_845_n572# a_853_n560# 0.07fF
C473 a_93_26# b1 0.13fF
C474 w_n114_n1393# a_n47_n1382# 0.08fF
C475 a_n169_n349# a_n105_n390# 0.16fF
C476 a_789_n2# a_852_174# 0.05fF
C477 a_14_139# a_99_201# 0.40fF
C478 w_162_n986# a_168_n1052# 0.19fF
C479 s2o gnd 0.23fF
C480 vddc2 a_517_n491# 2.46fF
C481 p1 a_673_n77# 0.05fF
C482 a_n99_n1099# vdd 0.78fF
C483 a_n3_n947# clk 0.05fF
C484 g1 g3 0.29fF
C485 b4 a4 0.49fF
C486 p2 p4 0.19fF
C487 w_775_n133# a_842_n122# 0.08fF
C488 a_14_139# gnd 0.24fF
C489 w_63_n1799# b4i 0.09fF
C490 a_739_n1491# a_802_n1315# 0.05fF
C491 a_517_n491# a_548_n492# 1.24fF
C492 vddc2 a_566_n630# 0.02fF
C493 b4 gnd 0.23fF
C494 w_n136_n610# clk 0.10fF
C495 clk m2_2_n1512# 0.03fF
C496 w_198_n821# p3 1.14fF
C497 vddc3 a_589_n837# 1.07fF
C498 w_1046_163# vdd 0.11fF
C499 w_196_n392# b2 0.31fF
C500 w_781_57# a_789_69# 0.07fF
C501 a_n76_n78# vdd 0.78fF
C502 a_890_n231# a_913_n297# 0.08fF
C503 w_1057_n133# a_1064_n230# 0.08fF
C504 a_940_66# gnd 0.21fF
C505 a_940_66# s1o 0.13fF
C506 w_504_n499# g1 0.08fF
C507 a_n99_n1194# clk 0.05fF
C508 a_548_n492# a_566_n630# 1.24fF
C509 b1 vdd11 0.03fF
C510 b4 a_69_n1617# 0.13fF
C511 c0 vdd 0.44fF
C512 a_330_117# gnd 0.24fF
C513 w_n105_n300# a_n182_n322# 0.08fF
C514 s3 p3 0.52fF
C515 c2 gndc2 0.24fF
C516 clk w_87_183# 0.10fF
C517 vdds1 a_673_n77# 0.45fF
C518 p1 a_516_n838# 0.08fF
C519 p2 p3 0.39fF
C520 a_n110_n1558# a_n110_n1487# 0.40fF
C521 g3 a_168_n1052# 0.17fF
C522 a_330_117# a_315_86# 0.21fF
C523 a_n210_n146# gnd 0.24fF
C524 p2 a_658_n289# 0.05fF
C525 a_1004_n563# gnd 0.21fF
C526 a_853_n631# a_913_n631# 0.08fF
C527 vdds3 a_734_n545# 0.45fF
C528 w_n132_n504# vdd 0.70fF
C529 w_493_n1362# a_543_n1355# 0.62fF
C530 a_n50_n1558# a_n5_n1557# 0.08fF
C531 w_n218_n87# a_n210_n146# 0.08fF
C532 a_153_n309# gnd1 0.71fF
C533 a_200_n1654# a_69_n1656# 0.08fF
C534 a_658_n289# gnds2 0.22fF
C535 a_739_n1491# clk 0.05fF
C536 w_n7_n341# a_n99_n215# 0.08fF
C537 a_529_n251# c1 0.07fF
C538 a_92_48# w_191_75# 0.17fF
C539 a_315_160# clk 0.05fF
C540 a_890_n1423# vdd 0.44fF
C541 a_n68_n669# clk 0.07fF
C542 w_735_n1326# a_850_n1424# 0.17fF
C543 a2 vdd 0.44fF
C544 w_n112_n783# a_n108_n948# 0.09fF
C545 w_n214_19# a_n147_30# 0.08fF
C546 b2 a_169_n461# 0.05fF
C547 a_n97_n1142# a_n99_n1194# 0.08fF
C548 a_506_n1632# a_525_n1632# 1.03fF
C549 a_506_n1355# a_543_n1355# 2.13fF
C550 a_172_n1419# gnd4 0.22fF
C551 a_43_n880# a3 0.13fF
C552 a_3_n881# a_n3_n947# 0.21fF
C553 a1i a_n210_n75# 0.05fF
C554 w_n105_n1259# b3i 0.09fF
C555 a_26_n880# vdd 0.78fF
C556 a_317_115# clk 0.07fF
C557 b1 w_191_75# 0.08fF
C558 g1 vdd1 0.44fF
C559 clk m2_236_n1660# 0.03fF
C560 a_951_n1058# clk 0.05fF
C561 w_n151_n81# clk 0.10fF
C562 w_1046_163# s1o 0.09fF
C563 a_29_96# clk 0.05fF
C564 a_884_n297# clk 0.05fF
C565 a_169_n890# gnd3 0.22fF
C566 vddc3 a_516_n838# 4.50fF
C567 a_24_n1490# a_24_n1557# 0.23fF
C568 c0 gnd 0.23fF
C569 w_n132_n504# a_n65_n493# 0.08fF
C570 w_n136_n610# a_n128_n669# 0.08fF
C571 a_n108_n948# gnd 0.24fF
C572 gndc2 a_529_n630# 0.78fF
C573 w_731_n1432# clk 0.10fF
C574 p2 g3 0.29fF
C575 b4 a_172_n1419# 0.05fF
C576 a_964_n564# a_958_n630# 0.21fF
C577 s4 a_725_n1062# 0.20fF
C578 w_500_n844# c0 0.06fF
C579 a_529_n251# a_512_n251# 0.41fF
C580 c1 gndc1 0.21fF
C581 w_n112_n783# a_26_n880# 0.17fF
C582 w_n111_n233# clk 0.10fF
C583 w_504_n499# p2 0.42fF
C584 a_779_n298# a_839_n298# 0.08fF
C585 w_201_n1350# b4 0.23fF
C586 w_849_n466# a_853_n560# 0.08fF
C587 clk m2_27_n900# 0.03fF
C588 a_900_65# a_894_n1# 0.21fF
C589 a_890_n1423# gnd 0.21fF
C590 a_957_n992# a_980_n991# 0.05fF
C591 a2 gnd 0.23fF
C592 w_735_n1326# vdd 0.70fF
C593 w_134_n112# b1 0.07fF
C594 a_913_n230# vdd 0.78fF
C595 clk m2_377_88# 0.03fF
C596 a_n99_n1194# a_n96_n1244# 0.40fF
C597 w_500_n844# c3 0.46fF
C598 a_n50_n1558# clk 0.07fF
C599 g1 p2 0.49fF
C600 a_23_n601# vdd 0.44fF
C601 a_n169_n349# clk 0.05fF
C602 a_n128_n669# a_n68_n669# 0.08fF
C603 a_900_65# vdd 0.41fF
C604 a_32_n1114# clk 0.05fF
C605 w_n51_n1493# a_n47_n1382# 0.07fF
C606 w_849_n466# s3o 0.08fF
C607 a_n76_n78# a_n59_n78# 0.18fF
C608 a_n105_n145# clk 0.05fF
C609 g4 gnd44 0.25fF
C610 w_n214_19# vdd 0.70fF
C611 a_26_n947# gnd 0.21fF
C612 a_105_134# vdd 0.44fF
C613 p3 b3 0.52fF
C614 a_906_n1059# a_951_n1058# 0.08fF
C615 a_n184_n277# a_n93_n282# 0.05fF
C616 gndc4 a_596_n1632# 0.55fF
C617 a_570_n1089# a_608_n1088# 0.82fF
C618 w_838_n233# clk 0.10fF
C619 a_n99_n79# a_n105_n145# 0.21fF
C620 clk m2_891_n252# 0.03fF
C621 w_n69_n604# a_n68_n669# 0.08fF
C622 w_842_n894# a_906_n1059# 0.09fF
C623 a_393_69# vdd 0.78fF
C624 w_838_n1000# a_846_n1059# 0.08fF
C625 gndc1 a_512_n251# 0.41fF
C626 a_964_n564# vdd 0.41fF
C627 a_850_n1424# a_873_n1423# 0.05fF
C628 w_735_n1326# c4 0.09fF
C629 a_n110_n1487# vdd 0.44fF
C630 a_171_n1581# a_178_n1581# 0.47fF
C631 c0 p1 0.83fF
C632 w_n114_n1393# a_n110_n1487# 0.08fF
C633 a_789_n2# w_785_163# 0.09fF
C634 vdd a_69_n1656# 0.41fF
C635 a_846_n1059# clk 0.05fF
C636 a_900_65# w_785_163# 0.17fF
C637 w_n105_n1259# a_n97_n1142# 0.09fF
C638 vdds4 a_725_n1062# 0.45fF
C639 a_930_n230# s2o 0.13fF
C640 a_739_n1491# a_739_n1420# 0.40fF
C641 w_162_n986# b3 0.06fF
C642 clk m2_70_n1143# 0.03fF
C643 a3i a_n108_n877# 0.05fF
C644 w_1124_n894# a_1131_n991# 0.08fF
C645 p4 a4 0.98fF
C646 a_n99_n1116# a_33_n1137# 0.21fF
C647 s1 a_789_69# 0.05fF
C648 a_n17_n602# a_n23_n668# 0.21fF
C649 vdd4 a_172_n1419# 0.45fF
C650 p1 a_147_n147# 0.20fF
C651 a_n184_n277# clk 0.05fF
C652 a_789_n2# gnd 0.24fF
C653 w_63_n1799# a_69_n1734# 0.09fF
C654 w_163_n1736# a_72_n1732# 0.07fF
C655 a_23_n601# gnd 0.21fF
C656 g2 a_168_n623# 0.17fF
C657 p1 a_512_n120# 0.09fF
C658 w_493_n1362# a_614_n1355# 0.56fF
C659 a_890_n231# a_884_n297# 0.21fF
C660 w_775_n133# s2o 0.08fF
C661 a_923_66# a_940_66# 0.18fF
C662 c0 g4 0.09fF
C663 w_493_n1362# a_506_n1355# 0.71fF
C664 a_394_47# vdd 0.44fF
C665 w_n7_n341# a_n184_n277# 0.09fF
C666 c3 s4 0.98fF
C667 a_561_n1632# a_596_n1632# 1.03fF
C668 a_873_n1423# vdd 0.78fF
C669 a_16_94# a_29_96# 0.08fF
C670 a_853_n631# a_853_n560# 0.40fF
C671 p3 a_734_n545# 0.05fF
C672 a_24_n1490# vdd 0.78fF
C673 w_731_n1432# a_739_n1420# 0.07fF
C674 w_912_n566# clk 0.10fF
C675 w_735_n1326# a_799_n1491# 0.09fF
C676 a_n169_n320# gnd 0.24fF
C677 w_n114_n1393# a_24_n1490# 0.17fF
C678 w_500_n844# p3 0.69fF
C679 a2 a_n105_n390# 0.13fF
C680 a_n97_n1142# a_n96_n1192# 0.40fF
C681 a_315_86# a_393_69# 0.05fF
C682 vddc1 c1 0.41fF
C683 a_512_n120# a_529_n251# 0.91fF
C684 w_n5_n1196# a_n96_n1192# 0.07fF
C685 w_n105_n1259# a_n96_n1244# 0.08fF
C686 a_725_n1062# gnds4 0.22fF
C687 a_987_n563# a_1004_n563# 0.18fF
C688 a_846_n1059# a_906_n1059# 0.08fF
C689 vddc3 c3 0.44fF
C690 clk m2_874_n1443# 0.03fF
C691 a_14_139# clk 0.05fF
C692 w_n151_n81# a_n150_n146# 0.08fF
C693 a_26_n880# a_43_n880# 0.18fF
C694 w_n132_n504# a_n128_n598# 0.08fF
C695 gnd b4i 0.12fF
C696 p1 p4 0.19fF
C697 a_909_n883# vdd 0.44fF
C698 w_848_63# clk 0.10fF
C699 a_43_n880# a_26_n947# 0.16fF
C700 g3 gnd33 0.25fF
C701 a3 a_169_n890# 0.05fF
C702 b3 vdd3 0.03fF
C703 a_330_117# clk 0.05fF
C704 w_63_n1799# vdd 0.70fF
C705 w_n214_19# a_n59_n78# 0.17fF
C706 b3 a_168_n1052# 0.42fF
C707 w_1046_163# a_1053_66# 0.08fF
C708 a_394_47# gnd 0.21fF
C709 p4 a_172_n1419# 0.20fF
C710 a_69_n1656# a_71_n1682# 0.05fF
C711 a_n210_n146# clk 0.05fF
C712 a_734_n545# gnds3 0.22fF
C713 a_n184_n277# a_n182_n322# 0.08fF
C714 w_493_n1362# g2 0.07fF
C715 a_14_65# a_29_67# 0.08fF
C716 w_504_n499# a_517_n491# 0.21fF
C717 p1 p3 0.38fF
C718 a_890_n1423# a_873_n1490# 0.16fF
C719 s4 p4 0.52fF
C720 w_n112_n783# a_n48_n948# 0.09fF
C721 w_500_n844# g3 0.08fF
C722 w_n116_n889# a_n108_n877# 0.07fF
C723 w_492_n126# p1 0.06fF
C724 a_1131_n991# vdd 0.44fF
C725 w_504_n499# a_566_n630# 0.35fF
C726 s1 a_673_n77# 0.20fF
C727 w_201_n1350# p4 1.14fF
C728 w_500_n844# a_608_n1088# 0.96fF
C729 a_779_n298# a_779_n227# 0.40fF
C730 a_n184_n351# clk 0.02fF
C731 a_33_n1137# gnd 0.24fF
C732 a_n76_n145# gnd 0.21fF
C733 p4 g4 0.09fF
C734 w_849_n466# a_1004_n563# 0.17fF
C735 clk m2_375_111# 0.03fF
C736 a_400_222# vdd 0.44fF
C737 a_n17_n602# vdd 0.41fF
C738 w_198_n821# b3 0.23fF
C739 a_n150_n146# a_n105_n145# 0.08fF
C740 a_779_n298# gnd 0.24fF
C741 a_n48_n948# gnd 0.23fF
C742 w_n7_n341# a_n184_n351# 0.17fF
C743 g1 gnd1 0.25fF
C744 a_852_174# vdd 0.44fF
C745 w_500_n844# g1 0.06fF
C746 w_492_n126# a_529_n251# 0.24fF
C747 p3 g4 0.09fF
C748 w_n114_n1393# a_n110_n1558# 0.09fF
C749 a_n99_n79# a_n76_n78# 0.05fF
C750 a_n108_n948# clk 0.05fF
C751 a_175_n623# gnd22 0.71fF
C752 a_406_155# vdd 0.44fF
C753 b2i gnd 0.12fF
C754 clk m2_901_44# 0.03fF
C755 w_842_n894# a_846_n988# 0.08fF
C756 a_14_65# vdd 0.41fF
C757 a_916_n455# vdd 0.44fF
C758 w_155_n858# a_169_n890# 0.08fF
C759 p2 a_552_n838# 0.08fF
C760 w_63_n1799# a_69_n1617# 0.17fF
C761 w_1124_n894# vdd 0.11fF
C762 clk m2_68_n1120# 0.03fF
C763 a_n50_n1558# a_1_n1491# 0.05fF
C764 a_n169_n349# a_n106_n368# 0.23fF
C765 a_14_139# w_191_75# 0.09fF
C766 p1 g3 0.29fF
C767 a_1131_n991# gnd 0.23fF
C768 a_852_174# w_785_163# 0.08fF
C769 a_913_n230# a_930_n230# 0.18fF
C770 p4 vdds4 0.03fF
C771 w_1_n1263# clk 0.10fF
C772 c0i a_400_222# 0.05fF
C773 w_504_n499# p1 0.08fF
C774 a_n59_n78# a_n76_n145# 0.16fF
C775 a1 b1 0.49fF
C776 a_n147_30# vdd 0.44fF
C777 w_842_n894# s4o 0.08fF
C778 a_1131_n563# vdd 0.44fF
C779 w_912_n566# a_913_n631# 0.08fF
C780 a_839_n298# gnd 0.23fF
C781 a_980_n991# a_980_n1058# 0.23fF
C782 w_63_n1799# a_71_n1682# 0.09fF
C783 w_n111_n233# a_n99_n215# 0.07fF
C784 a_315_160# a_317_115# 0.08fF
C785 a_24_n1557# gnd 0.21fF
C786 a_23_n601# a_6_n668# 0.16fF
C787 p1 g1 0.56fF
C788 w_781_57# a_789_n2# 0.08fF
C789 a_26_n947# clk 0.05fF
C790 w_n7_n341# a2 0.08fF
C791 a_n182_n322# a_n184_n351# 0.05fF
C792 w_905_n994# a_909_n883# 0.07fF
C793 a_850_n1424# vdd 0.41fF
C794 w_775_n133# a_913_n230# 0.17fF
C795 a_900_65# a_923_66# 0.05fF
C796 a_14_139# a_16_94# 0.08fF
C797 a_n23_n668# gnd 0.24fF
C798 w_735_n1326# a_802_n1315# 0.08fF
C799 w_731_n1432# a_739_n1491# 0.08fF
C800 g3 g4 0.09fF
C801 a_n110_n1558# gnd 0.24fF
C802 a_543_n1355# a_578_n1355# 2.06fF
C803 w_848_63# a_849_n2# 0.08fF
C804 w_n132_n504# b2 0.08fF
C805 gnd a_200_n1654# 0.21fF
C806 s3 gnd 0.12fF
C807 w_771_n239# a_779_n298# 0.08fF
C808 vdd11 a_147_n147# 0.45fF
C809 a_n99_n1116# vdd 0.41fF
C810 w_n105_n1259# a_n99_n1194# 0.09fF
C811 a_69_n1617# a_200_n1654# 0.16fF
C812 s3 a_734_n545# 0.20fF
C813 vddc3 a_608_n1088# 0.03fF
C814 clk w_388_204# 0.10fF
C815 clk m2_851_n1445# 0.03fF
C816 b2 a2 0.58fF
C817 w_n214_19# a1i 0.09fF
C818 w_500_n844# p2 0.53fF
C819 w_154_n425# vdd2 0.08fF
C820 a_147_n147# gnd11 0.22fF
C821 g1 a_529_n251# 0.19fF
C822 vddc1 a_512_n120# 1.80fF
C823 w_n132_n504# a_n128_n669# 0.09fF
C824 a_964_n564# a_987_n563# 0.05fF
C825 g1 g4 0.09fF
C826 a_846_n1059# a_846_n988# 0.40fF
C827 c1 s2 0.98fF
C828 a_789_n2# clk 0.05fF
C829 a_1131_n563# gnd 0.23fF
C830 gndc3 a_534_n1089# 0.70fF
C831 w_158_n1387# a_172_n1419# 0.08fF
C832 a_3_n881# a_26_n880# 0.05fF
C833 a_69_n1656# a_201_n1677# 0.21fF
C834 gnd a_69_n1734# 0.24fF
C835 a_900_65# clk 0.02fF
C836 w_n105_n1259# a_n99_n1077# 0.17fF
C837 a_3_n881# a_26_n947# 0.08fF
C838 a_n210_n146# a_n150_n146# 0.08fF
C839 b3 vdd 0.44fF
C840 s1 c0 0.98fF
C841 a_873_n1423# a_873_n1490# 0.23fF
C842 c4o a_1024_n1423# 0.13fF
C843 g2 a_529_n630# 0.23fF
C844 w_838_n233# a_842_n122# 0.07fF
C845 w_n114_n1393# vdd 0.70fF
C846 a_n99_n1077# a_32_n1114# 0.16fF
C847 w_n116_n889# a_n108_n948# 0.08fF
C848 w_n214_19# a_n99_n79# 0.17fF
C849 a_29_67# gnd 0.21fF
C850 a_n96_n1192# a_n99_n1194# 0.05fF
C851 w_162_n557# b2 0.06fF
C852 a_964_n564# clk 0.02fF
C853 a_958_n630# gnd 0.24fF
C854 a_n184_n277# a_n99_n215# 0.40fF
C855 a_n169_n320# clk 0.05fF
C856 g2 a_561_n1632# 0.08fF
C857 w_165_n1515# a_171_n1581# 0.19fF
C858 w_n132_n504# a_6_n601# 0.17fF
C859 a_69_n1656# clk 0.02fF
C860 w_1_n1263# a_n96_n1244# 0.07fF
C861 p1 p2 0.49fF
C862 g1 gndc1 0.05fF
C863 vddc4 c4 0.41fF
C864 w_176_n77# p1 1.92fF
C865 w_n118_n1499# a_n110_n1487# 0.07fF
C866 a_997_n991# vdd 0.44fF
C867 a_1004_n563# a_987_n630# 0.16fF
C868 gndc4 a_561_n1632# 0.71fF
C869 w_n112_n783# vdd 0.70fF
C870 vdd w_785_163# 0.70fF
C871 b2i a_n128_n598# 0.05fF
C872 b2 a_23_n601# 0.13fF
C873 a_71_n1682# a_69_n1734# 0.08fF
C874 a_799_n1491# a_850_n1424# 0.05fF
C875 a_779_n227# vdd 0.44fF
C876 a2 a_168_n623# 0.12fF
C877 w_165_n1515# a4 0.06fF
C878 w_849_n466# a_964_n564# 0.17fF
C879 a_168_n1052# a_175_n1052# 0.47fF
C880 a_894_n1# gnd 0.24fF
C881 a_940_66# a_923_n1# 0.16fF
C882 a_n65_n493# vdd 0.44fF
C883 gndc3 c3 0.21fF
C884 w_134_n112# a_147_n147# 0.07fF
C885 a_1064_n230# vdd 0.44fF
C886 w_842_n894# a_846_n1059# 0.09fF
C887 a_99_201# vdd 0.44fF
C888 a4 vdd 0.44fF
C889 w_492_n126# vddc1 0.44fF
C890 clk m2_981_n1011# 0.03fF
C891 w_n114_n1393# a4 0.08fF
C892 a_n184_n351# a_n106_n368# 0.05fF
C893 b3 gnd 0.23fF
C894 p2 g4 0.09fF
C895 s1o vdd 0.44fF
C896 w_n49_n883# a_n48_n948# 0.08fF
C897 w_775_n133# a_779_n298# 0.09fF
C898 w_1017_n1326# a_1024_n1423# 0.08fF
C899 p3 a_169_n890# 0.20fF
C900 a_315_86# vdd 0.41fF
C901 a_69_n1617# vdd 0.44fF
C902 w_493_n1362# a_578_n1355# 0.57fF
C903 a_14_139# w_87_183# 0.08fF
C904 a_315_160# w_492_96# 0.09fF
C905 w_500_n844# a_552_n838# 0.50fF
C906 a_33_n1137# clk 0.05fF
C907 a_997_n991# gnd 0.21fF
C908 w_1124_n466# s3o 0.09fF
C909 a4 a_171_n1581# 0.12fF
C910 a_n76_n145# clk 0.05fF
C911 w_162_n557# a_168_n623# 0.19fF
C912 a_890_n231# a_913_n230# 0.05fF
C913 w_493_n1362# c0 0.07fF
C914 a_578_n1355# a_614_n1355# 2.06fF
C915 w_n111_n233# a_n184_n277# 0.08fF
C916 s1o w_785_163# 0.08fF
C917 a_317_115# w_492_96# 0.09fF
C918 a_n99_n79# a_n76_n145# 0.08fF
C919 a_105_134# w_191_75# 0.08fF
C920 a_406_155# w_394_137# 0.07fF
C921 a_n182_n322# a_n169_n320# 0.08fF
C922 w_842_n894# a_980_n991# 0.17fF
C923 c4 gnd 0.12fF
C924 w_735_n1326# a_739_n1420# 0.08fF
C925 a_779_n298# clk 0.05fF
C926 a_6_n601# a_23_n601# 0.18fF
C927 a_24_n1490# a_41_n1490# 0.18fF
C928 a_n48_n948# clk 0.07fF
C929 c0i gnd 0.12fF
C930 a_789_n2# a_849_n2# 0.08fF
C931 w_140_n243# b1 0.06fF
C932 a_1064_n230# gnd 0.23fF
C933 a_n17_n602# a_6_n668# 0.08fF
C934 w_n105_n1259# a_n96_n1192# 0.08fF
C935 w_775_n133# a_839_n298# 0.09fF
C936 a_849_n2# a_900_65# 0.05fF
C937 vddc2 c2 0.41fF
C938 a_168_n623# vdd22 1.15fF
C939 a4 gnd 0.23fF
C940 clk m2_25_n1510# 0.03fF
C941 w_196_n392# a2 0.14fF
C942 a_n59_n78# vdd 0.44fF
C943 a_n108_n948# a_n45_n772# 0.05fF
C944 a_913_n230# a_913_n297# 0.23fF
C945 a_33_n1137# a_n97_n1142# 0.08fF
C946 s1o gnd 0.23fF
C947 g3 a_596_n1632# 0.08fF
C948 b1 a_147_n147# 0.05fF
C949 a_16_94# a_105_134# 0.40fF
C950 a_317_115# a_330_117# 0.08fF
C951 w_169_n1803# a_69_n1734# 0.08fF
C952 a_69_n1617# gnd 0.21fF
C953 clk w_93_116# 0.10fF
C954 vdds2 a_658_n289# 0.45fF
C955 gndc3 a_516_n1088# 0.82fF
C956 b1 a_146_n309# 0.42fF
C957 a_330_88# a_393_69# 0.23fF
C958 a_913_n631# a_964_n564# 0.05fF
C959 a_839_n298# clk 0.07fF
C960 w_165_n1515# g4 0.06fF
C961 a_799_n1491# gnd 0.23fF
C962 a_850_n1424# a_873_n1490# 0.08fF
C963 a_24_n1557# clk 0.05fF
C964 a_n17_n602# clk 0.02fF
C965 a_n99_n1077# a_n99_n1099# 0.18fF
C966 a_n105_n390# vdd 0.44fF
C967 w_n214_19# a_n150_n146# 0.09fF
C968 a2 a_169_n461# 0.05fF
C969 a_n48_n948# a_3_n881# 0.05fF
C970 gnd a_71_n1682# 0.23fF
C971 a_n23_n668# clk 0.05fF
C972 a_n110_n1558# clk 0.05fF
C973 clk m2_7_n621# 0.03fF
C974 a_200_n1654# clk 0.05fF
C975 w_1_n1263# a_n99_n1194# 0.08fF
C976 a_n210_n146# a_n210_n75# 0.40fF
C977 a_43_n880# vdd 0.44fF
C978 a_1004_n563# s3o 0.13fF
C979 w_771_n239# a_779_n227# 0.07fF
C980 a_909_n883# a_906_n1059# 0.40fF
C981 g2 gnd22 0.25fF
C982 vdd3 a_169_n890# 0.45fF
C983 w_n118_n1499# a_n110_n1558# 0.08fF
C984 a_14_65# clk 0.02fF
C985 w_493_n1362# p4 0.94fF
C986 a_n59_n78# gnd 0.21fF
C987 c0 g2 0.42fF
C988 p1 a_517_n491# 0.06fF
C989 vddc3 a_552_n838# 1.44fF
C990 a_41_n1490# a_24_n1557# 0.16fF
C991 w_n132_n504# a_n68_n669# 0.09fF
C992 a_957_n992# vdd 0.41fF
C993 g4 a_171_n1581# 0.17fF
C994 a4 a_172_n1419# 0.05fF
C995 p4 a_614_n1355# 0.08fF
C996 a_330_88# a_394_47# 0.16fF
C997 a_964_n564# a_987_n630# 0.08fF
C998 w_500_n844# p1 0.06fF
C999 a_n128_n598# vdd 0.44fF
C1000 w_n112_n783# a_43_n880# 0.17fF
C1001 gndc3 a_608_n1088# 0.21fF
C1002 w_493_n1362# p3 0.85fF
C1003 w_849_n466# s3 0.09fF
C1004 w_849_n466# a_916_n455# 0.08fF
C1005 a_n47_n1382# a_n50_n1558# 0.40fF
C1006 clk m2_958_n1013# 0.03fF
C1007 w_201_n1350# a4 0.13fF
C1008 s4 gnd 0.12fF
C1009 a_900_65# a_923_n1# 0.08fF
C1010 a_n184_n351# a_n169_n349# 0.08fF
C1011 a_72_n1784# b4i 0.05fF
C1012 a_69_n1734# clk 0.05fF
C1013 a_n105_n390# gnd 0.21fF
C1014 a_930_n230# vdd 0.44fF
C1015 clk m2_76_67# 0.03fF
C1016 p2 b2 0.56fF
C1017 w_n105_n1259# a_n99_n1099# 0.17fF
C1018 a_850_n1424# clk 0.02fF
C1019 a_633_n1632# c4 0.08fF
C1020 a2i gnd 0.12fF
C1021 a_29_67# clk 0.05fF
C1022 a_43_n880# gnd 0.21fF
C1023 a_958_n630# clk 0.05fF
C1024 a_n99_n1099# a_32_n1114# 0.23fF
C1025 a_923_66# vdd 0.78fF
C1026 s2 a_658_n289# 0.20fF
C1027 w_1017_n1326# c4o 0.09fF
C1028 a_n99_n1116# clk 0.02fF
C1029 a_1053_66# vdd 0.44fF
C1030 a_n93_n282# vdd 0.44fF
C1031 w_775_n133# vdd 0.70fF
C1032 a_29_67# a_93_26# 0.16fF
C1033 p2 a_543_n1355# 0.09fF
C1034 a_315_160# w_388_204# 0.08fF
C1035 a_987_n563# vdd 0.78fF
C1036 a_802_n1315# vdd 0.44fF
C1037 w_500_n844# vddc3 0.92fF
C1038 w_140_n243# a1 0.06fF
C1039 w_735_n1326# a_739_n1491# 0.09fF
C1040 a_175_n1052# gnd33 0.71fF
C1041 w_162_n557# g2 0.06fF
C1042 a_839_n298# a_890_n231# 0.05fF
C1043 a_n5_n1557# gnd 0.24fF
C1044 w_493_n1362# g3 0.07fF
* C1045 m2_238_n1683# Gnd 0.04fF **FLOATING
* C1046 m2_236_n1660# Gnd 0.04fF **FLOATING
* C1047 m2_874_n1443# Gnd 0.04fF **FLOATING
* C1048 m2_851_n1445# Gnd 0.04fF **FLOATING
* C1049 m2_25_n1510# Gnd 0.04fF **FLOATING
* C1050 m2_2_n1512# Gnd 0.04fF **FLOATING
* C1051 m2_70_n1143# Gnd 0.04fF **FLOATING
* C1052 m2_68_n1120# Gnd 0.04fF **FLOATING
* C1053 m2_981_n1011# Gnd 0.04fF **FLOATING
* C1054 m2_958_n1013# Gnd 0.04fF **FLOATING
* C1055 m2_27_n900# Gnd 0.04fF **FLOATING
* C1056 m2_4_n902# Gnd 0.04fF **FLOATING
* C1057 m2_988_n583# Gnd 0.04fF **FLOATING
* C1058 m2_965_n585# Gnd 0.04fF **FLOATING
* C1059 m2_7_n621# Gnd 0.04fF **FLOATING
* C1060 m2_n16_n623# Gnd 0.04fF **FLOATING
* C1061 m2_n122_n349# Gnd 0.04fF **FLOATING
* C1062 m2_n124_n326# Gnd 0.04fF **FLOATING
* C1063 m2_914_n250# Gnd 0.04fF **FLOATING
* C1064 m2_891_n252# Gnd 0.04fF **FLOATING
* C1065 m2_924_46# Gnd 0.04fF **FLOATING
* C1066 m2_901_44# Gnd 0.04fF **FLOATING
* C1067 m2_n75_n98# Gnd 0.04fF **FLOATING
* C1068 m2_n98_n100# Gnd 0.04fF **FLOATING
* C1069 m2_76_67# Gnd 0.04fF **FLOATING
* C1070 m2_377_88# Gnd 0.04fF **FLOATING
* C1071 m2_74_90# Gnd 0.04fF **FLOATING
* C1072 m2_375_111# Gnd 0.04fF **FLOATING
C1073 clk Gnd 9.90fF
C1074 b4i Gnd 1.02fF
C1075 a_72_n1784# Gnd 0.19fF
C1076 a_69_n1734# Gnd 1.78fF
C1077 a_72_n1732# Gnd 0.14fF
C1078 a_71_n1682# Gnd 1.64fF
C1079 a_201_n1677# Gnd 0.24fF
C1080 a_69_n1656# Gnd 1.45fF
C1081 a_200_n1654# Gnd 0.22fF
C1082 a_69_n1639# Gnd 0.84fF
C1083 gnd Gnd 30.21fF
C1084 a_873_n1490# Gnd 0.14fF
C1085 a_844_n1490# Gnd 0.24fF
C1086 a_1024_n1423# Gnd 0.37fF
C1087 vdd Gnd 19.52fF
C1088 c4o Gnd 1.15fF
C1089 a_890_n1423# Gnd 0.84fF
C1090 a_873_n1423# Gnd 0.84fF
C1091 a_850_n1424# Gnd 1.45fF
C1092 a_799_n1491# Gnd 1.64fF
C1093 a_802_n1315# Gnd 0.14fF
C1094 a_739_n1420# Gnd 0.19fF
C1095 a_739_n1491# Gnd 1.78fF
C1096 c4 Gnd 1.92fF
C1097 a_633_n1632# Gnd 2.61fF
C1098 a_596_n1632# Gnd 0.33fF
C1099 a_561_n1632# Gnd 0.33fF
C1100 a_578_n1355# Gnd 0.00fF
C1101 a_525_n1632# Gnd 0.35fF
C1102 a_506_n1632# Gnd 0.24fF
C1103 gndc4 Gnd 1.03fF
C1104 a_69_n1617# Gnd 0.84fF
C1105 gnd44 Gnd 0.54fF
C1106 a_178_n1581# Gnd 0.17fF
C1107 vdd44 Gnd 0.09fF
C1108 a_24_n1557# Gnd 0.22fF
C1109 a_171_n1581# Gnd 0.63fF
C1110 gnd4 Gnd 0.11fF
C1111 a_n5_n1557# Gnd 0.24fF
C1112 a_543_n1355# Gnd 0.03fF
C1113 a_506_n1355# Gnd 0.02fF
C1114 vddc4 Gnd 0.34fF
C1115 a_172_n1419# Gnd 0.51fF
C1116 vdd4 Gnd 0.04fF
C1117 a_41_n1490# Gnd 0.84fF
C1118 a_24_n1490# Gnd 0.84fF
C1119 a_1_n1491# Gnd 1.45fF
C1120 a_n50_n1558# Gnd 1.64fF
C1121 a_n47_n1382# Gnd 0.14fF
C1122 a_n110_n1487# Gnd 0.00fF
C1123 a_n110_n1558# Gnd 1.78fF
C1124 a4i Gnd 1.02fF
C1125 a4 Gnd 4.82fF
C1126 b4 Gnd 2.31fF
C1127 b3i Gnd 1.02fF
C1128 a_n96_n1244# Gnd 0.19fF
C1129 a_n99_n1194# Gnd 1.78fF
C1130 a_n96_n1192# Gnd 0.14fF
C1131 g4 Gnd 2.97fF
C1132 a_n97_n1142# Gnd 1.64fF
C1133 a_33_n1137# Gnd 0.24fF
C1134 a_n99_n1116# Gnd 1.45fF
C1135 a_32_n1114# Gnd 0.22fF
C1136 a_n99_n1099# Gnd 0.84fF
C1137 gnds4 Gnd 0.11fF
C1138 a_980_n1058# Gnd 0.22fF
C1139 a_951_n1058# Gnd 0.24fF
C1140 a_725_n1062# Gnd 0.59fF
C1141 vdds4 Gnd 0.12fF
C1142 p4 Gnd 13.05fF
C1143 a_1131_n991# Gnd 0.37fF
C1144 s4o Gnd 1.15fF
C1145 a_997_n991# Gnd 0.84fF
C1146 a_980_n991# Gnd 0.84fF
C1147 a_957_n992# Gnd 1.45fF
C1148 a_906_n1059# Gnd 1.64fF
C1149 a_909_n883# Gnd 0.14fF
C1150 a_846_n988# Gnd 0.19fF
C1151 a_846_n1059# Gnd 1.78fF
C1152 s4 Gnd 3.39fF
C1153 c3 Gnd 2.07fF
C1154 a_608_n1088# Gnd 2.16fF
C1155 a_570_n1089# Gnd 0.30fF
C1156 a_589_n837# Gnd 0.13fF
C1157 a_534_n1089# Gnd 0.30fF
C1158 a_516_n1088# Gnd 0.19fF
C1159 gndc3 Gnd 1.21fF
C1160 a_n99_n1077# Gnd 0.84fF
C1161 gnd33 Gnd 0.54fF
C1162 a_175_n1052# Gnd 0.17fF
C1163 vdd33 Gnd 0.09fF
C1164 a_168_n1052# Gnd 0.63fF
C1165 gnd3 Gnd 0.09fF
C1166 a_516_n838# Gnd 0.09fF
C1167 vddc3 Gnd 0.46fF
C1168 a_26_n947# Gnd 0.22fF
C1169 a_169_n890# Gnd 0.51fF
C1170 vdd3 Gnd 0.04fF
C1171 a_n3_n947# Gnd 0.24fF
C1172 b3 Gnd 2.68fF
C1173 a3 Gnd 4.78fF
C1174 a_43_n880# Gnd 0.84fF
C1175 a_26_n880# Gnd 0.84fF
C1176 a_3_n881# Gnd 1.45fF
C1177 a_n48_n948# Gnd 1.64fF
C1178 a_n45_n772# Gnd 0.14fF
C1179 a_n108_n877# Gnd 0.00fF
C1180 a_n108_n948# Gnd 1.78fF
C1181 a3i Gnd 1.03fF
C1182 g3 Gnd 6.23fF
C1183 a_987_n630# Gnd 0.22fF
C1184 a_958_n630# Gnd 0.24fF
C1185 a_529_n630# Gnd 0.27fF
C1186 gnd22 Gnd 0.54fF
C1187 a_175_n623# Gnd 0.17fF
C1188 gnds3 Gnd 0.11fF
C1189 a_1131_n563# Gnd 0.37fF
C1190 s3o Gnd 1.13fF
C1191 a_1004_n563# Gnd 0.84fF
C1192 a_987_n563# Gnd 0.84fF
C1193 a_964_n564# Gnd 1.45fF
C1194 a_913_n631# Gnd 1.64fF
C1195 a_916_n455# Gnd 0.14fF
C1196 a_853_n560# Gnd 0.19fF
C1197 a_734_n545# Gnd 0.59fF
C1198 vdds3 Gnd 0.12fF
C1199 gndc2 Gnd 1.70fF
C1200 p3 Gnd 17.26fF
C1201 a_853_n631# Gnd 1.78fF
C1202 s3 Gnd 3.39fF
C1203 c2 Gnd 1.43fF
C1204 a_566_n630# Gnd 0.85fF
C1205 a_6_n668# Gnd 0.14fF
C1206 vdd22 Gnd 0.09fF
C1207 a_168_n623# Gnd 0.63fF
C1208 a_n23_n668# Gnd 0.16fF
C1209 g2 Gnd 7.47fF
C1210 vddc2 Gnd 0.44fF
C1211 gnd2 Gnd 0.09fF
C1212 a_23_n601# Gnd 0.84fF
C1213 a_6_n601# Gnd 0.84fF
C1214 a_n17_n602# Gnd 1.45fF
C1215 a_n68_n669# Gnd 1.64fF
C1216 a_n65_n493# Gnd 0.14fF
C1217 a_n128_n598# Gnd 0.19fF
C1218 a_n128_n669# Gnd 1.78fF
C1219 b2i Gnd 1.01fF
C1220 a_169_n461# Gnd 0.52fF
C1221 vdd2 Gnd 0.04fF
C1222 a_n105_n390# Gnd 0.84fF
C1223 a2 Gnd 6.24fF
C1224 b2 Gnd 2.18fF
C1225 a_n106_n368# Gnd 0.84fF
C1226 a_n169_n349# Gnd 0.22fF
C1227 a_n184_n351# Gnd 1.45fF
C1228 a_n169_n320# Gnd 0.24fF
C1229 a_913_n297# Gnd 0.22fF
C1230 gnds2 Gnd 0.11fF
C1231 a_884_n297# Gnd 0.24fF
C1232 gnd1 Gnd 0.54fF
C1233 a_153_n309# Gnd 0.17fF
C1234 a_n93_n282# Gnd 0.14fF
C1235 a_658_n289# Gnd 0.59fF
C1236 vdds2 Gnd 0.12fF
C1237 p2 Gnd 10.05fF
C1238 a_1064_n230# Gnd 0.37fF
C1239 s2o Gnd 1.15fF
C1240 a_930_n230# Gnd 0.84fF
C1241 a_913_n230# Gnd 0.84fF
C1242 a_890_n231# Gnd 1.45fF
C1243 a_839_n298# Gnd 1.64fF
C1244 a_842_n122# Gnd 0.14fF
C1245 a_779_n227# Gnd 0.19fF
C1246 a_512_n251# Gnd 0.10fF
C1247 gndc1 Gnd 0.64fF
C1248 a_n182_n322# Gnd 1.64fF
C1249 vdd1 Gnd 0.09fF
C1250 a_n99_n215# Gnd 0.19fF
C1251 a_n184_n277# Gnd 1.78fF
C1252 a2i Gnd 1.01fF
C1253 a_146_n309# Gnd 0.63fF
C1254 gnd11 Gnd 0.11fF
C1255 a_779_n298# Gnd 1.78fF
C1256 s2 Gnd 3.39fF
C1257 gnds1 Gnd 0.10fF
C1258 c1 Gnd 1.94fF
C1259 a_529_n251# Gnd 1.41fF
C1260 a_512_n120# Gnd 0.06fF
C1261 vddc1 Gnd 0.24fF
C1262 g1 Gnd 8.11fF
C1263 a_923_n1# Gnd 0.22fF
C1264 a_894_n1# Gnd 0.24fF
C1265 a_673_n77# Gnd 0.59fF
C1266 vdds1 Gnd 0.12fF
C1267 a_147_n147# Gnd 0.52fF
C1268 vdd11 Gnd 0.03fF
C1269 a_n76_n145# Gnd 0.22fF
C1270 b1 Gnd 2.05fF
C1271 a_n105_n145# Gnd 0.24fF
C1272 p1 Gnd 12.10fF
C1273 c0 Gnd 8.93fF
C1274 a_93_26# Gnd 0.84fF
C1275 a_394_47# Gnd 0.84fF
C1276 a_92_48# Gnd 0.84fF
C1277 a_29_67# Gnd 0.22fF
C1278 a1 Gnd 5.09fF
C1279 a_n59_n78# Gnd 0.84fF
C1280 a_n76_n78# Gnd 0.84fF
C1281 a_n99_n79# Gnd 1.45fF
C1282 a_n150_n146# Gnd 1.64fF
C1283 a_n147_30# Gnd 0.14fF
C1284 a_n210_n75# Gnd 0.00fF
C1285 a_n210_n146# Gnd 1.78fF
C1286 a1i Gnd 1.01fF
C1287 a_393_69# Gnd 0.84fF
C1288 a_330_88# Gnd 0.22fF
C1289 a_14_65# Gnd 1.45fF
C1290 a_29_96# Gnd 0.24fF
C1291 a_315_86# Gnd 1.45fF
C1292 a_330_117# Gnd 0.24fF
C1293 a_1053_66# Gnd 0.37fF
C1294 a_105_134# Gnd 0.14fF
C1295 a_16_94# Gnd 1.64fF
C1296 a_406_155# Gnd 0.14fF
C1297 a_317_115# Gnd 1.64fF
C1298 s1o Gnd 1.08fF
C1299 a_940_66# Gnd 0.84fF
C1300 a_923_66# Gnd 0.84fF
C1301 a_900_65# Gnd 1.45fF
C1302 a_849_n2# Gnd 1.64fF
C1303 a_852_174# Gnd 0.14fF
C1304 a_789_69# Gnd 0.19fF
C1305 a_99_201# Gnd 0.19fF
C1306 a_14_139# Gnd 1.78fF
C1307 b1i Gnd 1.01fF
C1308 a_789_n2# Gnd 1.78fF
C1309 s1 Gnd 3.38fF
C1310 a_400_222# Gnd 0.19fF
C1311 a_315_160# Gnd 1.78fF
C1312 c0i Gnd 1.04fF
C1313 w_169_n1803# Gnd 1.87fF
C1314 w_163_n1736# Gnd 1.87fF
C1315 w_63_n1799# Gnd 12.07fF
C1316 w_165_n1515# Gnd 4.60fF
C1317 w_n51_n1493# Gnd 0.13fF
C1318 w_n118_n1499# Gnd 0.87fF
C1319 w_798_n1426# Gnd 1.87fF
C1320 w_731_n1432# Gnd 1.87fF
C1321 w_1017_n1326# Gnd 1.81fF
C1322 w_735_n1326# Gnd 12.07fF
C1323 w_158_n1387# Gnd 1.52fF
C1324 w_n114_n1393# Gnd 12.07fF
C1325 w_201_n1350# Gnd 3.15fF
C1326 w_1_n1263# Gnd 1.87fF
C1327 w_n5_n1196# Gnd 1.87fF
C1328 w_493_n1362# Gnd 45.34fF
C1329 w_n105_n1259# Gnd 12.07fF
C1330 w_905_n994# Gnd 1.87fF
C1331 w_838_n1000# Gnd 0.01fF
C1332 w_162_n986# Gnd 4.60fF
C1333 w_1124_n894# Gnd 1.81fF
C1334 w_842_n894# Gnd 12.07fF
C1335 w_500_n844# Gnd 34.45fF
C1336 w_155_n858# Gnd 1.52fF
C1337 w_n49_n883# Gnd 0.20fF
C1338 w_n116_n889# Gnd 1.21fF
C1339 w_198_n821# Gnd 3.15fF
C1340 w_n112_n783# Gnd 12.07fF
C1341 w_912_n566# Gnd 1.87fF
C1342 w_845_n572# Gnd 1.87fF
C1343 w_162_n557# Gnd 4.60fF
C1344 w_n69_n604# Gnd 1.87fF
C1345 w_n136_n610# Gnd 1.87fF
C1346 w_1124_n466# Gnd 1.81fF
C1347 w_n132_n504# Gnd 12.07fF
C1348 w_849_n466# Gnd 12.07fF
C1349 w_504_n499# Gnd 19.38fF
C1350 w_196_n392# Gnd 4.22fF
C1351 w_154_n425# Gnd 1.41fF
C1352 w_838_n233# Gnd 1.87fF
C1353 w_771_n239# Gnd 1.87fF
C1354 w_140_n243# Gnd 4.60fF
C1355 w_n7_n341# Gnd 12.07fF
C1356 w_n105_n300# Gnd 1.87fF
C1357 w_n111_n233# Gnd 1.87fF
C1358 w_1057_n133# Gnd 1.81fF
C1359 w_775_n133# Gnd 12.07fF
C1360 w_492_n126# Gnd 10.46fF
C1361 w_134_n112# Gnd 0.69fF
C1362 w_176_n77# Gnd 4.76fF
C1363 w_n151_n81# Gnd 0.13fF
C1364 w_n218_n87# Gnd 0.84fF
C1365 w_848_63# Gnd 1.87fF
C1366 w_781_57# Gnd 1.87fF
C1367 w_n214_19# Gnd 12.07fF
C1368 w_1046_163# Gnd 1.81fF
C1369 w_785_163# Gnd 12.07fF
C1370 w_492_96# Gnd 12.07fF
C1371 w_394_137# Gnd 1.87fF
C1372 w_388_204# Gnd 1.87fF
C1373 w_191_75# Gnd 12.07fF
C1374 w_93_116# Gnd 1.87fF
C1375 w_87_183# Gnd 1.87fF

.tran 0.1n 50n
* .measure tran delays0 TRIG v(b1) VAL=0.9 RISE=1 TARG v(s4) VAL=0.9 rise=1
* .measure tran delays1 TRIG v(b2) VAL=0.9 RISE=1 TARG v(s2) VAL=0.9 RISE=1
* .measure tran delays2 TRIG v(b3) VAL=0.9 RISE=1 TARG v(s3) VAL=0.9 RISE=1
* .measure tran delays3 TRIG v(b4) VAL=0.9 RISE=1 TARG v(s4) VAL=0.9 RISE=1
* .measure tran carry4 TRIG v(c0) VAL=0.9 RISE=3 TARG v(c4) VAL=0.9 RISE=1

.control
set hcopypscolor=1
set color0=white
set color1=black
run

set curplottitle="Sanjana Sheela - 20231012027- postlayout"
* plot v(a1i) v(a2i)+2 v(a3i)+4 v(a4i)+6 v(clk)+8
* plot v(b1i) v(b2i)+2 v(b3i)+4 v(b4i)+6 v(clk)+8 v(c0i)-2
* plot v(a1) v(a2)+2 v(a3)+4 v(a4)+6 v(clk)+8
* plot v(b1) v(b2)+2 v(b3)+4 v(b4)+6 v(clk)+8 v(c0)-2
* plot v(s1o) v(s2o)+2 v(s3o)+4 v(s4o)+6 v(c4o)+8 v(clk)+10
* plot v(g1) v(p1)+2 v(g2)+4 v(p2)+6 v(g3)+8 v(p3)+10 v(g4)+12 v(p4)+14
* plot v(c0)-2 v(c1) v(c2)+2 v(c3)+4 v(c4)+6
plot v(s1) v(s2)+2 v(s3)+4 v(s4)+6 

* plot v(a1i) v(a1)+2 v(clk)+4
* plot v(a2i) v(a2)+2 v(clk)+4
* plot v(a3i) v(a3)+2 v(clk)+4
* plot v(a4i) v(a4)+2 v(clk)+4

* plot v(b1i) v(b1)+2 v(clk)+4
* plot v(b2i) v(b2)+2 v(clk)+4
* plot v(b3i) v(b3)+2 v(clk)+4
* plot v(b4i) v(b4)+2 v(clk)+4

* plot v(c0i) v(c0)+2 v(clk)+4

* plot v(s1) v(s1o)+2 v(clk)+4
* plot v(s2) v(s2o)+2 v(clk)+4
* plot v(s3) v(s3o)+2 v(clk)+4
* plot v(s4) v(s4o)+2 v(clk)+4

* plot v(a1) v(b1)+2 v(p1)+4 
* plot v(a2) v(b2)+2 v(p2)+4 
* plot v(a3) v(b3)+2 v(p3)+4 
* plot v(a4) v(b4)+2 v(p4)+4

* plot v(a1) v(b1)+2 v(g1)+4 
* plot v(a2) v(b2)+2 v(g2)+4 
* plot v(a3) v(b3)+2 v(g3)+4 
* plot v(a4) v(b4)+2 v(g4)+4

* plot v(p1) v(g1)+2 v(c0)+4 v(c1)+6
* plot v(p2) v(g2)+2 v(c1)+4 v(c2)+6
* plot v(p3) v(g3)+2 v(c2)+4 v(c3)+6
* plot v(p4) v(g4)+2 v(c3)+4 v(c4)+6


* plot v(a1) v(b1)+2 v(c0)+4 v(p1)+6 v(g1)+8 v(s1)+10 v(c1)+12
* plot v(a2) v(b2)+2 v(c1)+4 v(p2)+6 v(g2)+8 v(s2)+10 v(c2)+12
* plot v(a3) v(b3)+2 v(c2)+4 v(p3)+6 v(g3)+8 v(s3)+10 v(c3)+12
* plot v(a4) v(b4)+2 v(c3)+4 v(p4)+6 v(g4)+8 v(s4)+10 v(c4)+12
.endc
.end

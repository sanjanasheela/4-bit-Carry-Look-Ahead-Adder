* Propagate and Generate Block
.include TSMC_180nm.txt

.param LAMBDA=0.09u
.param SUPPLY=1.8
.param width=1.8u
.param Wp = 2*width
.param Wn = width
.global gnd vdd

Vdd vdd gnd 'SUPPLY'
Va1 a1 gnd pulse(0 1.8 2n 0 0 2n 4n)
Va2 a2 gnd pulse(0 1.8 2n 0 0 4n 8n)
Va3 a3 gnd pulse(0 1.8 2n 0 0 8n 16n)
Va4 a4 gnd pulse(0 1.8 2n 0 0 16n 32n)

Vb1 b1 gnd pulse(0 1.8 2n 0 0 16n 32n)
Vb2 b2 gnd pulse(0 1.8 2n 0 0 8n 16n)
Vb3 b3 gnd pulse(0 1.8 2n 0 0 4n 8n)
Vb4 b4 gnd pulse(0 1.8 2n 0 0 2n 4n)

* SPICE3 file created from pgblock.ext - technology: scmos

.option scale=0.09u

M1000 gnd a_127_n743# g2 Gnd CMOSN w=20 l=2
+  ad=1580 pd=752 as=100 ps=50
M1001 p2 a2 b2 Vdd CMOSP w=40 l=2
+  ad=400 pd=180 as=200 ps=90
M1002 p3 b3 a3 Vdd CMOSP w=40 l=2
+  ad=400 pd=180 as=200 ps=90
M1003 p4 a4 a_121_n1415# Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=190 ps=96
M1004 a_120_n1577# a4 vdd w_114_n1511# CMOSP w=40 l=2
+  ad=400 pd=180 as=3200 ps=1440
M1005 g1 a_139_n309# vdd w_133_n243# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1006 a_140_n147# b1 vdd Vdd CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1007 a_146_n309# a1 a_139_n309# Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=200 ps=90
M1008 p3 a3 a_128_n1021# Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=190 ps=96
M1009 p4 b4 a4 Vdd CMOSP w=40 l=2
+  ad=400 pd=180 as=200 ps=90
M1010 a_120_n1577# b4 vdd w_114_n1511# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 gnd a_120_n1577# g4 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1012 gnd b2 a_134_n743# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1013 a_121_n1415# b4 gnd Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=0 ps=0
M1014 a_139_n309# b1 vdd w_133_n243# CMOSP w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1015 a_128_n1021# b3 vdd Vdd CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1016 a_134_n1183# a3 a_127_n1183# Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=200 ps=90
M1017 p1 a_140_n147# a1 Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=95 ps=48
M1018 g3 a_127_n1183# vdd w_121_n1117# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1019 p4 a_121_n1415# a4 Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=95 ps=48
M1020 gnd b3 a_134_n1183# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1021 gnd a_139_n309# g1 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1022 p2 b2 a2 Vdd CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1023 g2 a_127_n743# vdd w_121_n677# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1024 a_134_n743# a2 a_127_n743# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1025 p1 a1 b1 Vdd CMOSP w=40 l=2
+  ad=400 pd=180 as=200 ps=90
M1026 a_139_n309# a1 vdd w_133_n243# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 p2 a2 a_128_n581# Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=190 ps=96
M1028 p3 a_128_n1021# a3 Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=95 ps=48
M1029 p1 b1 a1 Vdd CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1030 a_140_n147# b1 gnd Gnd CMOSN w=19 l=2
+  ad=190 pd=96 as=0 ps=0
M1031 a_127_n743# b2 vdd w_121_n677# CMOSP w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1032 a_127_n1577# a4 a_120_n1577# Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=200 ps=90
M1033 p3 a3 b3 Vdd CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1034 g4 a_120_n1577# vdd w_114_n1511# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1035 a_128_n581# b2 vdd Vdd CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1036 gnd b4 a_127_n1577# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 a_121_n1415# b4 vdd Vdd CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1038 a_127_n1183# a3 vdd w_121_n1117# CMOSP w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1039 a_127_n743# a2 vdd w_121_n677# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1040 a_127_n1183# b3 vdd w_121_n1117# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 p4 a4 b4 Vdd CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1042 p2 a_128_n581# a2 Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=95 ps=48
M1043 a_128_n581# b2 gnd Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 gnd a_127_n1183# g3 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1045 p1 a1 a_140_n147# Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 gnd b1 a_146_n309# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1047 a_128_n1021# b3 gnd Gnd CMOSN w=19 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_114_n1511# vdd 0.39fF
C1 a2 a_128_n581# 0.05fF
C2 b2 p2 0.52fF
C3 w_121_n1117# b3 0.06fF
C4 a_128_n1021# vdd 0.45fF
C5 g2 gnd 0.25fF
C6 a_140_n147# p1 0.20fF
C7 a_121_n1415# vdd 0.45fF
C8 a_134_n1183# gnd 0.71fF
C9 w_114_n1511# g4 0.06fF
C10 g4 gnd 0.25fF
C11 b2 a_127_n743# 0.42fF
C12 a2 p2 0.98fF
C13 w_121_n1117# a3 0.06fF
C14 a_134_n743# gnd 0.71fF
C15 b2 vdd 0.03fF
C16 a_140_n147# gnd 0.22fF
C17 a_127_n1577# gnd 0.71fF
C18 b3 a3 0.49fF
C19 a_128_n581# p2 0.20fF
C20 a2 a_127_n743# 0.12fF
C21 a_139_n309# g1 0.17fF
C22 w_121_n677# b2 0.06fF
C23 b4 a4 0.49fF
C24 a2 vdd 0.02fF
C25 w_114_n1511# b4 0.06fF
C26 b3 a_128_n1021# 0.05fF
C27 a_127_n1183# g3 0.17fF
C28 a_139_n309# a_146_n309# 0.47fF
C29 w_121_n677# a2 0.06fF
C30 b4 a_121_n1415# 0.05fF
C31 a_128_n581# vdd 0.45fF
C32 a_127_n1183# vdd 1.15fF
C33 g1 gnd 0.25fF
C34 w_114_n1511# a4 0.06fF
C35 a_120_n1577# vdd 1.15fF
C36 a3 a_128_n1021# 0.05fF
C37 a_127_n1183# a_134_n1183# 0.47fF
C38 a4 a_121_n1415# 0.05fF
C39 a_128_n1021# gnd 0.22fF
C40 a_146_n309# gnd 0.71fF
C41 a_121_n1415# gnd 0.22fF
C42 a_120_n1577# g4 0.17fF
C43 b3 p3 0.52fF
C44 w_121_n1117# a_127_n1183# 0.19fF
C45 a_127_n743# vdd 1.15fF
C46 b4 p4 0.52fF
C47 g3 vdd 0.44fF
C48 w_133_n243# b1 0.06fF
C49 a_120_n1577# a_127_n1577# 0.47fF
C50 b1 vdd 0.03fF
C51 w_133_n243# vdd 0.39fF
C52 a3 p3 0.98fF
C53 b3 a_127_n1183# 0.42fF
C54 a_127_n743# g2 0.17fF
C55 w_121_n677# a_127_n743# 0.19fF
C56 g2 vdd 0.44fF
C57 a4 p4 0.98fF
C58 b4 a_120_n1577# 0.42fF
C59 b1 a1 0.49fF
C60 w_133_n243# a1 0.06fF
C61 a1 vdd 0.02fF
C62 w_121_n677# vdd 0.39fF
C63 vdd g4 0.44fF
C64 a_128_n1021# p3 0.20fF
C65 a3 a_127_n1183# 0.12fF
C66 a_127_n743# a_134_n743# 0.47fF
C67 w_121_n677# g2 0.06fF
C68 w_121_n1117# g3 0.06fF
C69 a_121_n1415# p4 0.20fF
C70 a4 a_120_n1577# 0.12fF
C71 a_128_n581# gnd 0.22fF
C72 b1 a_140_n147# 0.05fF
C73 a_140_n147# vdd 0.45fF
C74 w_114_n1511# a_120_n1577# 0.19fF
C75 w_121_n1117# vdd 0.39fF
C76 b2 a2 0.49fF
C77 b3 vdd 0.03fF
C78 b1 a_139_n309# 0.42fF
C79 w_133_n243# a_139_n309# 0.19fF
C80 a_139_n309# vdd 1.15fF
C81 a1 a_140_n147# 0.05fF
C82 b1 p1 0.52fF
C83 b4 vdd 0.03fF
C84 b2 a_128_n581# 0.05fF
C85 a3 vdd 0.02fF
C86 a1 a_139_n309# 0.12fF
C87 w_133_n243# g1 0.06fF
C88 g1 vdd 0.44fF
C89 a1 p1 0.98fF
C90 g3 gnd 0.25fF
C91 a4 vdd 0.02fF
C92 gnd Gnd 2.56fF
C93 a_127_n1577# Gnd 0.17fF
C94 g4 Gnd 0.31fF
C95 vdd Gnd 0.78fF
C96 a_120_n1577# Gnd 0.63fF
C97 p4 Gnd 2.52fF
C98 a_121_n1415# Gnd 0.59fF
C99 a4 Gnd 4.50fF
C100 b4 Gnd 2.06fF
C101 a_134_n1183# Gnd 0.17fF
C102 g3 Gnd 0.31fF
C103 a_127_n1183# Gnd 0.63fF
C104 p3 Gnd 2.52fF
C105 a_128_n1021# Gnd 0.59fF
C106 a3 Gnd 4.50fF
C107 b3 Gnd 2.06fF
C108 a_134_n743# Gnd 0.17fF
C109 g2 Gnd 0.31fF
C110 a_127_n743# Gnd 0.63fF
C111 p2 Gnd 2.52fF
C112 a2 Gnd 4.50fF
C113 b2 Gnd 0.20fF
C114 a_146_n309# Gnd 0.17fF
C115 g1 Gnd 0.31fF
C116 a_139_n309# Gnd 0.63fF
C117 p1 Gnd 2.52fF
C118 a_140_n147# Gnd 0.07fF
C119 a1 Gnd 4.50fF
C120 b1 Gnd 0.20fF
C121 w_114_n1511# Gnd 4.60fF
C122 w_121_n1117# Gnd 4.60fF
C123 w_121_n677# Gnd 4.60fF
C124 w_133_n243# Gnd 4.60fF
.tran 0.1n 40n

.control

run
set curplottitle="Sanjana Sheela - 20231012027- postlayout"
plot v(a1) v(b1)+2 v(p1)+4
plot v(a2) v(b2)+2 v(p2)+4
plot v(a3) v(b3)+2 v(p3)+4
plot v(a4) v(b4)+2 v(p4)+4

plot v(a1) v(b1)+2 v(g1)+4
plot v(a2) v(b2)+2 v(g2)+4
plot v(a3) v(b3)+2 v(g3)+4
plot v(a4) v(b4)+2 v(g4)+4

.endc
.end

.include TSMC_180nm.txt


.param LAMBDA=0.09u
.param SUPPLY=1.8
.param width=1.8u
.param Wp = 2*width
.param Wn = width
.global gnd vdd

Vdd vdd gnd 'SUPPLY'
Va1 p1 gnd pulse(0 1.8 2n 0 0 2n 4n)
Va2 p2 gnd pulse(0 1.8 2n 0 0 4n 8n)
Va3 p3 gnd pulse(0 1.8 2n 0 0 8n 16n)
Va4 p4 gnd pulse(0 1.8 2n 0 0 16n 32n)

Vb1 c1 gnd pulse(0 1.8 2n 0 0 16n 32n)
Vb2 c2 gnd pulse(0 1.8 2n 0 0 8n 16n)
Vb3 c3 gnd pulse(0 1.8 2n 0 0 4n 8n)
Vb4 c0 gnd pulse(0 1.8 2n 0 0 2n 4n)


.subckt inv X Y vdd gnd Wp Wn LAMBDA
M1 Y X vdd vdd CMOSP W={Wp} L={2*LAMBDA} 
+AS={5*Wp*LAMBDA} PS={10*LAMBDA+2*Wp} 
+AD={5*Wp*LAMBDA} PD={10*LAMBDA+2*Wp}
M2 Y X gnd gnd CMOSN W={Wn} L={2*LAMBDA} 
+AS={5*Wn*LAMBDA} PS={10*LAMBDA+2*Wn} 
+AD={5*Wn*LAMBDA} PD={10*LAMBDA+2*Wn}
.ends


.subckt xor y a b vdd gnd
X1 b b_bar vdd gnd wp wn LAMBDA inv
M1 y b a vdd CMOSP W={Wp} L={2*LAMBDA} 
+AS={5*Wp*LAMBDA} PS={10*LAMBDA+2*Wp} 
+AD={5*Wp*LAMBDA} PD={10*LAMBDA+2*Wp}
M2 y b_bar a gnd CMOSN W={Wn} L={2*LAMBDA} 
+AS={5*Wn*LAMBDA} PS={10*LAMBDA+2*Wn} 
+AD={5*Wn*LAMBDA} PD={10*LAMBDA+2*Wn}
M3 y a b vdd CMOSP W={Wp} L={2*LAMBDA} 
+AS={5*Wp*LAMBDA} PS={10*LAMBDA+2*Wp} 
+AD={5*Wp*LAMBDA} PD={10*LAMBDA+2*Wp}
M4 y a b_bar gnd CMOSN W={Wn} L={2*LAMBDA} 
+AS={5*Wn*LAMBDA} PS={10*LAMBDA+2*Wn} 
+AD={5*Wn*LAMBDA} PD={10*LAMBDA+2*Wn}
.ends


X1 s1 p1 c0 vdd gnd xor
X2 s2 p2 c1 vdd gnd xor
X3 s3 p3 c2 vdd gnd xor
X4 s4 p4 c3 vdd gnd xor

.tran 0.1n 32n

.control

runset curplottitle="Sanjana Sheela - 20231012027- prelayout"


plot v(c0) v(c1)+2 v(c2)+4 (c3)+6 
plot v(p1) v(p2)+2 v(p3)+4 (p4)+6 
plot v(s1) v(s2)+2 v(s3)+4 (s4)+6 

.endc
.end


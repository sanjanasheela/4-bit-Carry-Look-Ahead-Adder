magic
tech scmos
timestamp 1732094920
<< nwell >>
rect 724 -32 737 -31
rect 644 -100 766 -32
rect 644 -126 725 -100
rect 626 -565 775 -564
rect 626 -636 810 -565
rect 626 -700 721 -636
rect 545 -1187 741 -1012
rect 538 -1715 746 -1700
rect 538 -1918 745 -1715
<< ntransistor >>
rect 662 -251 664 -211
rect 679 -251 681 -211
rect 710 -250 712 -230
rect 752 -247 754 -227
rect 790 -680 792 -660
rect 637 -831 639 -771
rect 649 -831 651 -771
rect 668 -801 670 -771
rect 686 -831 688 -771
rect 705 -791 707 -771
rect 559 -1431 561 -1351
rect 577 -1432 579 -1352
rect 595 -1431 597 -1391
rect 613 -1432 615 -1352
rect 632 -1431 634 -1405
rect 651 -1431 653 -1351
rect 669 -1431 671 -1411
rect 702 -1431 704 -1411
rect 549 -2188 551 -2088
rect 568 -2188 570 -2088
rect 586 -2188 588 -2138
rect 604 -2188 606 -2088
rect 621 -2188 623 -2155
rect 639 -2188 641 -2088
rect 657 -2188 659 -2163
rect 676 -2188 678 -2088
rect 695 -2188 697 -2168
rect 731 -2188 733 -2168
<< ptransistor >>
rect 662 -120 664 -40
rect 679 -120 681 -40
rect 710 -120 712 -40
rect 752 -82 754 -42
rect 637 -692 639 -572
rect 649 -692 651 -572
rect 668 -693 670 -573
rect 686 -633 688 -573
rect 705 -693 707 -573
rect 790 -624 792 -584
rect 559 -1181 561 -1021
rect 577 -1181 579 -1021
rect 595 -1181 597 -1021
rect 613 -1101 615 -1021
rect 632 -1180 634 -1020
rect 651 -1074 653 -1020
rect 669 -1179 671 -1019
rect 702 -1060 704 -1020
rect 549 -1911 551 -1711
rect 568 -1911 570 -1711
rect 586 -1911 588 -1711
rect 604 -1811 606 -1711
rect 621 -1911 623 -1711
rect 639 -1777 641 -1711
rect 657 -1911 659 -1711
rect 676 -1761 678 -1711
rect 695 -1911 697 -1711
rect 731 -1765 733 -1725
<< ndiffusion >>
rect 661 -251 662 -211
rect 664 -251 665 -211
rect 678 -251 679 -211
rect 681 -251 682 -211
rect 709 -250 710 -230
rect 712 -250 713 -230
rect 751 -247 752 -227
rect 754 -247 755 -227
rect 789 -680 790 -660
rect 792 -680 793 -660
rect 636 -831 637 -771
rect 639 -831 649 -771
rect 651 -831 652 -771
rect 667 -801 668 -771
rect 670 -801 671 -771
rect 685 -831 686 -771
rect 688 -831 689 -771
rect 704 -791 705 -771
rect 707 -791 708 -771
rect 558 -1431 559 -1351
rect 561 -1431 562 -1351
rect 576 -1432 577 -1352
rect 579 -1432 580 -1352
rect 594 -1431 595 -1391
rect 597 -1431 598 -1391
rect 612 -1432 613 -1352
rect 615 -1432 616 -1352
rect 631 -1431 632 -1405
rect 634 -1431 635 -1405
rect 650 -1431 651 -1351
rect 653 -1431 654 -1351
rect 668 -1431 669 -1411
rect 671 -1431 672 -1411
rect 701 -1431 702 -1411
rect 704 -1431 705 -1411
rect 548 -2188 549 -2088
rect 551 -2188 552 -2088
rect 567 -2188 568 -2088
rect 570 -2188 571 -2088
rect 585 -2188 586 -2138
rect 588 -2188 589 -2138
rect 603 -2188 604 -2088
rect 606 -2188 607 -2088
rect 620 -2188 621 -2155
rect 623 -2188 624 -2155
rect 638 -2188 639 -2088
rect 641 -2188 642 -2088
rect 656 -2188 657 -2163
rect 659 -2188 660 -2163
rect 675 -2188 676 -2088
rect 678 -2188 679 -2088
rect 694 -2188 695 -2168
rect 697 -2188 698 -2168
rect 730 -2188 731 -2168
rect 733 -2188 734 -2168
<< pdiffusion >>
rect 661 -120 662 -40
rect 664 -120 665 -40
rect 678 -120 679 -40
rect 681 -120 682 -40
rect 709 -120 710 -40
rect 712 -120 713 -40
rect 751 -82 752 -42
rect 754 -82 755 -42
rect 636 -692 637 -572
rect 639 -692 642 -572
rect 646 -692 649 -572
rect 651 -692 652 -572
rect 667 -693 668 -573
rect 670 -693 671 -573
rect 685 -633 686 -573
rect 688 -633 689 -573
rect 704 -693 705 -573
rect 707 -693 708 -573
rect 789 -624 790 -584
rect 792 -624 793 -584
rect 558 -1181 559 -1021
rect 561 -1181 562 -1021
rect 576 -1181 577 -1021
rect 579 -1181 580 -1021
rect 594 -1181 595 -1021
rect 597 -1181 598 -1021
rect 612 -1101 613 -1021
rect 615 -1101 616 -1021
rect 631 -1180 632 -1020
rect 634 -1180 635 -1020
rect 650 -1074 651 -1020
rect 653 -1074 654 -1020
rect 668 -1179 669 -1019
rect 671 -1179 672 -1019
rect 701 -1060 702 -1020
rect 704 -1060 705 -1020
rect 548 -1911 549 -1711
rect 551 -1911 552 -1711
rect 567 -1911 568 -1711
rect 570 -1911 571 -1711
rect 585 -1911 586 -1711
rect 588 -1911 589 -1711
rect 603 -1811 604 -1711
rect 606 -1811 607 -1711
rect 620 -1911 621 -1711
rect 623 -1911 624 -1711
rect 638 -1777 639 -1711
rect 641 -1777 642 -1711
rect 656 -1911 657 -1711
rect 659 -1911 660 -1711
rect 675 -1761 676 -1711
rect 678 -1761 679 -1711
rect 694 -1911 695 -1711
rect 697 -1911 698 -1711
rect 730 -1765 731 -1725
rect 733 -1765 734 -1725
<< ndcontact >>
rect 657 -251 661 -211
rect 665 -251 669 -211
rect 674 -251 678 -211
rect 682 -251 686 -211
rect 705 -250 709 -230
rect 713 -250 717 -230
rect 747 -247 751 -227
rect 755 -247 759 -227
rect 785 -680 789 -660
rect 793 -680 797 -660
rect 632 -831 636 -771
rect 652 -831 656 -771
rect 663 -801 667 -771
rect 671 -801 675 -771
rect 681 -831 685 -771
rect 689 -831 693 -771
rect 700 -791 704 -771
rect 708 -791 712 -771
rect 554 -1431 558 -1351
rect 562 -1431 566 -1351
rect 572 -1432 576 -1352
rect 580 -1432 584 -1352
rect 590 -1431 594 -1391
rect 598 -1431 602 -1391
rect 608 -1432 612 -1352
rect 616 -1432 620 -1352
rect 627 -1431 631 -1405
rect 635 -1431 639 -1405
rect 646 -1431 650 -1351
rect 654 -1431 658 -1351
rect 664 -1431 668 -1411
rect 672 -1431 676 -1411
rect 697 -1431 701 -1411
rect 705 -1431 709 -1411
rect 544 -2188 548 -2088
rect 552 -2188 556 -2088
rect 563 -2188 567 -2088
rect 571 -2188 575 -2088
rect 581 -2188 585 -2138
rect 589 -2188 593 -2138
rect 599 -2188 603 -2088
rect 607 -2188 611 -2088
rect 616 -2188 620 -2155
rect 624 -2188 628 -2155
rect 634 -2188 638 -2088
rect 642 -2188 646 -2088
rect 652 -2188 656 -2163
rect 660 -2188 664 -2163
rect 671 -2188 675 -2088
rect 679 -2188 683 -2088
rect 690 -2188 694 -2168
rect 698 -2188 702 -2168
rect 726 -2188 730 -2168
rect 734 -2188 738 -2168
<< pdcontact >>
rect 657 -120 661 -40
rect 665 -120 669 -40
rect 674 -120 678 -40
rect 682 -120 686 -40
rect 705 -120 709 -40
rect 713 -120 717 -40
rect 747 -82 751 -42
rect 755 -82 759 -42
rect 632 -692 636 -572
rect 642 -692 646 -572
rect 652 -692 656 -572
rect 663 -693 667 -573
rect 671 -693 675 -573
rect 681 -633 685 -573
rect 689 -633 693 -573
rect 700 -693 704 -573
rect 708 -693 712 -573
rect 785 -624 789 -584
rect 793 -624 797 -584
rect 554 -1181 558 -1021
rect 562 -1181 566 -1021
rect 572 -1181 576 -1021
rect 580 -1181 584 -1021
rect 590 -1181 594 -1021
rect 598 -1181 602 -1021
rect 608 -1101 612 -1021
rect 616 -1101 620 -1021
rect 627 -1180 631 -1020
rect 635 -1180 639 -1020
rect 646 -1074 650 -1020
rect 654 -1074 658 -1020
rect 664 -1179 668 -1019
rect 672 -1179 676 -1019
rect 697 -1060 701 -1020
rect 705 -1060 709 -1020
rect 544 -1911 548 -1711
rect 552 -1911 556 -1711
rect 563 -1911 567 -1711
rect 571 -1911 575 -1711
rect 581 -1911 585 -1711
rect 589 -1911 593 -1711
rect 599 -1811 603 -1711
rect 607 -1811 611 -1711
rect 616 -1911 620 -1711
rect 624 -1911 628 -1711
rect 634 -1777 638 -1711
rect 642 -1777 646 -1711
rect 652 -1911 656 -1711
rect 660 -1911 664 -1711
rect 671 -1761 675 -1711
rect 679 -1761 683 -1711
rect 690 -1911 694 -1711
rect 698 -1911 702 -1711
rect 726 -1765 730 -1725
rect 734 -1765 738 -1725
<< polysilicon >>
rect 662 -40 664 -37
rect 679 -40 681 -37
rect 710 -40 712 -37
rect 752 -42 754 -39
rect 662 -211 664 -120
rect 679 -211 681 -120
rect 710 -230 712 -120
rect 752 -227 754 -82
rect 662 -254 664 -251
rect 679 -254 681 -251
rect 710 -253 712 -250
rect 752 -252 754 -247
rect 637 -572 639 -569
rect 649 -572 651 -569
rect 668 -573 670 -569
rect 686 -573 688 -570
rect 705 -573 707 -570
rect 637 -771 639 -692
rect 649 -771 651 -692
rect 790 -584 792 -569
rect 790 -660 792 -624
rect 790 -683 792 -680
rect 668 -771 670 -693
rect 686 -771 688 -693
rect 705 -771 707 -693
rect 668 -805 670 -801
rect 705 -795 707 -791
rect 637 -834 639 -831
rect 649 -834 651 -831
rect 686 -834 688 -831
rect 559 -1021 561 -1018
rect 577 -1021 579 -1018
rect 595 -1021 597 -1018
rect 613 -1021 615 -1018
rect 632 -1020 634 -1017
rect 651 -1020 653 -1017
rect 669 -1019 671 -1016
rect 559 -1351 561 -1181
rect 577 -1352 579 -1181
rect 559 -1434 561 -1431
rect 595 -1391 597 -1181
rect 613 -1352 615 -1101
rect 577 -1435 579 -1432
rect 595 -1435 597 -1431
rect 632 -1405 634 -1180
rect 651 -1351 653 -1074
rect 702 -1020 704 -1017
rect 669 -1411 671 -1179
rect 702 -1411 704 -1060
rect 613 -1435 615 -1432
rect 632 -1434 634 -1431
rect 651 -1435 653 -1431
rect 669 -1435 671 -1431
rect 702 -1434 704 -1431
rect 549 -1711 551 -1708
rect 568 -1711 570 -1707
rect 586 -1711 588 -1707
rect 604 -1711 606 -1707
rect 621 -1711 623 -1708
rect 639 -1711 641 -1707
rect 657 -1711 659 -1708
rect 676 -1711 678 -1708
rect 695 -1711 697 -1708
rect 549 -2088 551 -1911
rect 568 -2088 570 -1911
rect 586 -2138 588 -1911
rect 604 -2088 606 -1811
rect 621 -2155 623 -1911
rect 639 -2088 641 -1777
rect 657 -2163 659 -1911
rect 676 -2088 678 -1761
rect 731 -1725 733 -1722
rect 695 -2168 697 -1911
rect 731 -2168 733 -1765
rect 549 -2191 551 -2188
rect 568 -2191 570 -2188
rect 586 -2191 588 -2188
rect 604 -2191 606 -2188
rect 621 -2191 623 -2188
rect 639 -2191 641 -2188
rect 657 -2191 659 -2188
rect 676 -2191 678 -2188
rect 695 -2191 697 -2188
rect 731 -2191 733 -2188
<< polycontact >>
rect 658 -137 662 -133
rect 675 -175 679 -171
rect 706 -208 710 -204
rect 748 -172 752 -167
rect 633 -708 637 -704
rect 645 -721 649 -717
rect 782 -651 790 -645
rect 664 -735 668 -731
rect 682 -749 686 -745
rect 701 -760 705 -756
rect 554 -1198 559 -1191
rect 572 -1217 577 -1210
rect 590 -1235 595 -1228
rect 608 -1256 613 -1249
rect 627 -1278 632 -1271
rect 646 -1305 651 -1298
rect 664 -1334 669 -1327
rect 698 -1309 702 -1305
rect 544 -1955 549 -1950
rect 563 -1969 568 -1964
rect 581 -1986 586 -1981
rect 599 -2000 604 -1995
rect 616 -2016 621 -2011
rect 634 -2029 639 -2024
rect 652 -2046 657 -2041
rect 671 -2060 676 -2055
rect 690 -2076 695 -2071
rect 726 -1965 731 -1959
<< polypplus >>
rect 686 -693 688 -633
<< metal1 >>
rect 644 -33 766 -29
rect 657 -40 661 -33
rect 682 -40 686 -33
rect 451 -81 455 -80
rect 237 -86 455 -81
rect 451 -171 455 -86
rect 669 -45 674 -40
rect 674 -123 678 -120
rect 705 -123 709 -120
rect 674 -128 709 -123
rect 747 -42 751 -33
rect 520 -137 658 -133
rect 713 -167 717 -120
rect 755 -131 759 -82
rect 755 -135 787 -131
rect 451 -175 486 -171
rect 493 -175 675 -171
rect 713 -172 748 -167
rect 522 -208 706 -204
rect 237 -248 451 -244
rect 522 -244 527 -208
rect 457 -248 527 -244
rect 669 -216 674 -211
rect 713 -221 717 -172
rect 705 -225 717 -221
rect 705 -230 709 -225
rect 755 -227 759 -135
rect 686 -250 705 -246
rect 657 -266 661 -251
rect 713 -266 717 -250
rect 747 -266 751 -247
rect 644 -270 764 -266
rect 626 -566 810 -560
rect 632 -572 636 -566
rect 652 -572 656 -566
rect 308 -593 312 -592
rect 284 -598 312 -593
rect 308 -745 312 -598
rect 689 -573 693 -566
rect 642 -695 646 -692
rect 675 -577 681 -573
rect 681 -641 685 -633
rect 675 -645 700 -641
rect 785 -584 789 -566
rect 793 -645 797 -624
rect 712 -651 782 -645
rect 793 -651 829 -645
rect 793 -660 797 -651
rect 785 -685 789 -680
rect 663 -695 666 -693
rect 642 -698 666 -695
rect 521 -708 633 -704
rect 493 -721 645 -717
rect 458 -735 664 -731
rect 307 -749 426 -745
rect 432 -749 682 -745
rect 284 -760 400 -756
rect 408 -760 701 -756
rect 708 -764 712 -693
rect 663 -768 685 -764
rect 663 -771 667 -768
rect 681 -771 685 -768
rect 700 -768 712 -764
rect 733 -691 812 -685
rect 700 -771 704 -768
rect 656 -775 663 -771
rect 632 -839 636 -831
rect 671 -839 675 -801
rect 693 -775 700 -771
rect 708 -839 712 -791
rect 733 -839 737 -691
rect 624 -845 737 -839
rect 545 -1014 741 -1008
rect 554 -1021 558 -1014
rect 580 -1021 584 -1014
rect 616 -1021 620 -1014
rect 654 -1020 658 -1014
rect 308 -1167 312 -1166
rect 279 -1172 312 -1167
rect 307 -1298 312 -1172
rect 566 -1026 572 -1021
rect 602 -1025 608 -1021
rect 608 -1107 612 -1101
rect 608 -1111 627 -1107
rect 639 -1025 646 -1020
rect 646 -1085 650 -1074
rect 646 -1089 664 -1085
rect 572 -1191 576 -1181
rect 590 -1191 594 -1181
rect 520 -1198 554 -1191
rect 571 -1195 594 -1191
rect 635 -1192 639 -1180
rect 664 -1192 668 -1179
rect 635 -1196 668 -1192
rect 697 -1020 701 -1014
rect 493 -1217 572 -1210
rect 458 -1235 590 -1228
rect 432 -1256 608 -1249
rect 408 -1278 627 -1271
rect 307 -1305 371 -1298
rect 378 -1305 646 -1298
rect 672 -1305 676 -1179
rect 705 -1305 709 -1060
rect 672 -1309 698 -1305
rect 705 -1309 789 -1305
rect 510 -1330 664 -1327
rect 279 -1334 664 -1330
rect 672 -1351 676 -1309
rect 566 -1431 572 -1426
rect 554 -1449 558 -1431
rect 584 -1356 608 -1352
rect 584 -1431 590 -1427
rect 584 -1432 594 -1431
rect 598 -1449 602 -1431
rect 620 -1356 646 -1352
rect 620 -1431 627 -1427
rect 658 -1355 678 -1351
rect 705 -1411 709 -1309
rect 658 -1431 664 -1427
rect 635 -1449 639 -1431
rect 672 -1449 676 -1431
rect 697 -1449 701 -1431
rect 531 -1455 714 -1449
rect 538 -1702 745 -1698
rect 544 -1711 548 -1702
rect 571 -1711 575 -1702
rect 607 -1711 611 -1702
rect 642 -1711 646 -1702
rect 679 -1711 683 -1702
rect 556 -1715 563 -1711
rect 556 -1910 563 -1907
rect 563 -1914 567 -1911
rect 581 -1914 585 -1911
rect 563 -1918 585 -1914
rect 593 -1715 599 -1711
rect 589 -1913 593 -1911
rect 628 -1715 634 -1711
rect 628 -1911 652 -1907
rect 664 -1716 671 -1711
rect 664 -1911 690 -1907
rect 726 -1725 730 -1702
rect 616 -1913 620 -1911
rect 589 -1918 620 -1913
rect 520 -1955 544 -1950
rect 698 -1958 702 -1911
rect 734 -1956 738 -1765
rect 698 -1959 725 -1958
rect 492 -1969 563 -1964
rect 698 -1965 726 -1959
rect 734 -1960 761 -1956
rect 457 -1986 581 -1981
rect 431 -2000 599 -1995
rect 407 -2016 616 -2011
rect 377 -2029 634 -2024
rect 344 -2046 652 -2041
rect 291 -2055 519 -2054
rect 291 -2060 671 -2055
rect 291 -2061 549 -2060
rect 500 -2072 690 -2071
rect 291 -2076 690 -2072
rect 544 -2193 548 -2188
rect 556 -2188 563 -2186
rect 575 -2093 599 -2088
rect 575 -2188 581 -2184
rect 611 -2092 634 -2088
rect 611 -2188 616 -2184
rect 646 -2092 671 -2088
rect 646 -2188 652 -2184
rect 698 -2154 702 -1965
rect 690 -2157 702 -2154
rect 690 -2168 694 -2157
rect 734 -2168 738 -1960
rect 683 -2188 690 -2184
rect 552 -2190 567 -2188
rect 589 -2193 593 -2188
rect 624 -2193 628 -2188
rect 660 -2193 664 -2188
rect 698 -2193 702 -2188
rect 726 -2193 730 -2188
rect 533 -2197 739 -2193
<< m123contact >>
rect 515 -137 520 -132
rect 486 -176 493 -170
rect 451 -249 457 -243
rect 514 -709 521 -703
rect 486 -722 493 -716
rect 451 -736 458 -730
rect 426 -749 432 -744
rect 400 -761 408 -756
rect 514 -1198 520 -1191
rect 487 -1217 493 -1210
rect 452 -1235 458 -1228
rect 426 -1256 432 -1249
rect 401 -1278 408 -1271
rect 371 -1305 378 -1298
rect 515 -1955 520 -1950
rect 487 -1969 492 -1964
rect 452 -1986 457 -1981
rect 426 -2000 431 -1995
rect 401 -2016 407 -2011
rect 371 -2029 377 -2024
rect 339 -2046 344 -2041
<< metal3 >>
rect 47 20 519 24
rect 515 -132 519 20
rect 452 -730 457 -249
rect 487 -716 492 -176
rect 515 -703 520 -137
rect 401 -1271 408 -761
rect 426 -1249 432 -749
rect 452 -1228 457 -736
rect 487 -1210 492 -722
rect 515 -1191 520 -709
rect 339 -2041 344 -1330
rect 371 -2024 377 -1305
rect 401 -2011 407 -1278
rect 426 -1995 431 -1256
rect 452 -1981 457 -1235
rect 487 -1964 492 -1217
rect 515 -1950 520 -1198
<< labels >>
rlabel metal3 100 22 104 23 5 c0
rlabel metal1 766 -134 770 -132 1 c1
rlabel metal1 822 -648 825 -647 1 c2
rlabel metal1 690 -269 690 -269 1 gndc1
rlabel metal1 679 -31 684 -29 1 vddc1
rlabel metal1 639 -843 642 -842 1 gndc2
rlabel metal1 675 -562 679 -561 1 vddc2
rlabel metal1 522 -1303 528 -1300 1 p3
rlabel metal1 727 -1307 735 -1305 1 c3
rlabel metal1 523 -1332 529 -1329 1 g3
rlabel metal1 588 -1011 596 -1010 1 vddc3
rlabel metal1 625 -1453 627 -1452 1 gndc3
rlabel metal1 520 -2059 521 -2058 1 p4
rlabel metal1 521 -2075 522 -2074 1 g4
rlabel metal1 745 -1958 745 -1958 1 c4
rlabel metal1 667 -1699 667 -1699 1 vddc4
rlabel metal1 611 -2196 611 -2196 1 gndc4
rlabel metal1 606 -759 616 -758 1 GG
rlabel metal1 396 -748 406 -746 1 p2
rlabel metal1 239 -246 239 -246 1 g1
rlabel metal1 247 -84 251 -83 1 p1
<< end >>

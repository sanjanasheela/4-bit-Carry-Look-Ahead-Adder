magic
tech scmos
timestamp 1732097814
<< ntransistor >>
rect 0 433 2 452
rect 30 433 32 452
rect -44 399 -42 418
rect 0 260 2 279
rect 30 260 32 279
rect -44 226 -42 245
rect -2 82 0 101
rect 28 82 30 101
rect -46 48 -44 67
rect -3 -73 -1 -54
rect 27 -73 29 -54
rect -47 -107 -45 -88
<< ptransistor >>
rect -44 441 -42 481
rect 0 475 2 515
rect 30 475 32 515
rect -44 268 -42 308
rect 0 302 2 342
rect 30 302 32 342
rect -46 90 -44 130
rect -2 124 0 164
rect 28 124 30 164
rect -47 -65 -45 -25
rect -3 -31 -1 9
rect 27 -31 29 9
<< ndiffusion >>
rect -1 433 0 452
rect 2 433 3 452
rect 29 433 30 452
rect 32 433 33 452
rect -45 399 -44 418
rect -42 399 -41 418
rect -1 260 0 279
rect 2 260 3 279
rect 29 260 30 279
rect 32 260 33 279
rect -45 226 -44 245
rect -42 226 -41 245
rect -3 82 -2 101
rect 0 82 1 101
rect 27 82 28 101
rect 30 82 31 101
rect -47 48 -46 67
rect -44 48 -43 67
rect -4 -73 -3 -54
rect -1 -73 0 -54
rect 26 -73 27 -54
rect 29 -73 30 -54
rect -48 -107 -47 -88
rect -45 -107 -44 -88
<< pdiffusion >>
rect -45 441 -44 481
rect -42 441 -41 481
rect -1 475 0 515
rect 2 475 3 515
rect 29 475 30 515
rect 32 475 33 515
rect -45 268 -44 308
rect -42 268 -41 308
rect -1 302 0 342
rect 2 302 3 342
rect 29 302 30 342
rect 32 302 33 342
rect -47 90 -46 130
rect -44 90 -43 130
rect -3 124 -2 164
rect 0 124 1 164
rect 27 124 28 164
rect 30 124 31 164
rect -48 -65 -47 -25
rect -45 -65 -44 -25
rect -4 -31 -3 9
rect -1 -31 0 9
rect 26 -31 27 9
rect 29 -31 30 9
<< ndcontact >>
rect -5 433 -1 452
rect 3 433 7 452
rect 25 433 29 452
rect 33 433 37 452
rect -49 399 -45 418
rect -41 399 -37 418
rect -5 260 -1 279
rect 3 260 7 279
rect 25 260 29 279
rect 33 260 37 279
rect -49 226 -45 245
rect -41 226 -37 245
rect -7 82 -3 101
rect 1 82 5 101
rect 23 82 27 101
rect 31 82 35 101
rect -51 48 -47 67
rect -43 48 -39 67
rect -8 -73 -4 -54
rect 0 -73 4 -54
rect 22 -73 26 -54
rect 30 -73 34 -54
rect -52 -107 -48 -88
rect -44 -107 -40 -88
<< pdcontact >>
rect -49 441 -45 481
rect -41 441 -37 481
rect -5 475 -1 515
rect 3 475 7 515
rect 25 475 29 515
rect 33 475 37 515
rect -49 268 -45 308
rect -41 268 -37 308
rect -5 302 -1 342
rect 3 302 7 342
rect 25 302 29 342
rect 33 302 37 342
rect -51 90 -47 130
rect -43 90 -39 130
rect -7 124 -3 164
rect 1 124 5 164
rect 23 124 27 164
rect 31 124 35 164
rect -52 -65 -48 -25
rect -44 -65 -40 -25
rect -8 -31 -4 9
rect 0 -31 4 9
rect 22 -31 26 9
rect 30 -31 34 9
<< polysilicon >>
rect 0 515 2 522
rect 30 515 32 518
rect -44 481 -42 484
rect 0 472 2 475
rect 0 452 2 455
rect 30 452 32 475
rect -44 418 -42 441
rect 0 426 2 433
rect 30 429 32 433
rect -44 395 -42 399
rect 0 342 2 349
rect 30 342 32 345
rect -44 308 -42 311
rect 0 299 2 302
rect 0 279 2 282
rect 30 279 32 302
rect -44 245 -42 268
rect 0 253 2 260
rect 30 256 32 260
rect -44 222 -42 226
rect -2 164 0 171
rect 28 164 30 167
rect -46 130 -44 133
rect -2 121 0 124
rect -2 101 0 104
rect 28 101 30 124
rect -46 67 -44 90
rect -2 75 0 82
rect 28 78 30 82
rect -46 44 -44 48
rect -3 9 -1 16
rect 27 9 29 12
rect -47 -25 -45 -22
rect -3 -34 -1 -31
rect -3 -54 -1 -51
rect 27 -54 29 -31
rect -47 -88 -45 -65
rect -3 -80 -1 -73
rect 27 -77 29 -73
rect -47 -111 -45 -107
<< polycontact >>
rect -4 518 0 522
rect 26 460 30 464
rect -48 426 -44 430
rect -4 426 0 430
rect -4 345 0 349
rect 26 287 30 291
rect -48 253 -44 257
rect -4 253 0 257
rect -6 167 -2 171
rect 24 109 28 113
rect -50 75 -46 79
rect -6 75 -2 79
rect -7 12 -3 16
rect 23 -46 27 -42
rect -51 -80 -47 -76
rect -7 -80 -3 -76
<< metal1 >>
rect -24 525 29 530
rect -24 522 -19 525
rect -63 518 -4 522
rect -63 430 -58 518
rect 25 515 29 525
rect -52 486 -35 490
rect -49 481 -45 486
rect -24 464 -19 495
rect -5 464 -1 475
rect 3 474 7 475
rect 33 465 37 475
rect -24 460 26 464
rect 33 460 42 465
rect 47 460 71 465
rect -41 430 -37 441
rect -5 452 -1 460
rect 33 452 37 460
rect -86 426 -48 430
rect -41 426 -4 430
rect -41 418 -37 426
rect -17 423 -13 426
rect 25 423 29 433
rect -17 418 29 423
rect -49 393 -45 399
rect -54 389 -35 393
rect -24 352 29 357
rect -24 349 -19 352
rect -63 345 -4 349
rect -63 257 -58 345
rect 25 342 29 352
rect -52 313 -35 317
rect -49 308 -45 313
rect -24 291 -19 322
rect -5 291 -1 302
rect 3 301 7 302
rect 33 292 37 302
rect -24 287 26 291
rect 33 287 42 292
rect 47 287 71 292
rect -41 257 -37 268
rect -5 279 -1 287
rect 33 279 37 287
rect -86 253 -48 257
rect -41 253 -4 257
rect -41 245 -37 253
rect -17 250 -13 253
rect 25 250 29 260
rect -17 245 29 250
rect -49 220 -45 226
rect -54 216 -35 220
rect -26 174 27 179
rect -26 171 -21 174
rect -65 167 -6 171
rect -65 79 -60 167
rect 23 164 27 174
rect -54 135 -37 139
rect -51 130 -47 135
rect -26 113 -21 144
rect -7 113 -3 124
rect 1 123 5 124
rect 31 114 35 124
rect -26 109 24 113
rect 31 109 40 114
rect 45 109 69 114
rect -43 79 -39 90
rect -7 101 -3 109
rect 31 101 35 109
rect -88 75 -50 79
rect -43 75 -6 79
rect -43 67 -39 75
rect -19 72 -15 75
rect 23 72 27 82
rect -19 67 27 72
rect -51 42 -47 48
rect -56 38 -37 42
rect -27 19 26 24
rect -27 16 -22 19
rect -66 12 -7 16
rect -66 -76 -61 12
rect 22 9 26 19
rect -55 -20 -38 -16
rect -52 -25 -48 -20
rect -27 -42 -22 -11
rect -8 -42 -4 -31
rect 0 -32 4 -31
rect 30 -41 34 -31
rect -27 -46 23 -42
rect 30 -46 39 -41
rect 44 -46 68 -41
rect -44 -76 -40 -65
rect -8 -54 -4 -46
rect 30 -54 34 -46
rect -89 -80 -51 -76
rect -44 -80 -7 -76
rect -44 -88 -40 -80
rect -20 -83 -16 -80
rect 22 -83 26 -73
rect -20 -88 26 -83
rect -52 -113 -48 -107
rect -57 -117 -38 -113
<< metal2 >>
rect 13 533 47 537
rect -88 495 -24 500
rect 13 474 18 533
rect 43 529 47 533
rect 8 469 18 474
rect 3 457 8 469
rect 42 465 47 529
rect 13 360 47 364
rect -88 322 -24 327
rect 13 301 18 360
rect 43 356 47 360
rect 8 296 18 301
rect 3 284 8 296
rect 42 292 47 356
rect 11 182 45 186
rect -90 144 -26 149
rect 11 123 16 182
rect 41 178 45 182
rect 6 118 16 123
rect 1 106 6 118
rect 40 114 45 178
rect 10 27 44 31
rect -91 -11 -27 -6
rect 10 -32 15 27
rect 40 23 44 27
rect 5 -37 15 -32
rect 0 -49 5 -37
rect 39 -41 44 23
<< m123contact >>
rect -24 495 -19 500
rect 3 469 8 474
rect 42 460 47 465
rect 3 452 8 457
rect -24 322 -19 327
rect 3 296 8 301
rect 42 287 47 292
rect 3 279 8 284
rect -26 144 -21 149
rect 1 118 6 123
rect 40 109 45 114
rect 1 101 6 106
rect -27 -11 -22 -6
rect 0 -37 5 -32
rect 39 -46 44 -41
rect 0 -54 5 -49
<< labels >>
rlabel metal1 -82 428 -82 428 1 c0
rlabel metal2 -83 497 -83 497 3 p1
rlabel metal1 -42 487 -42 487 1 vdd
rlabel metal1 -43 391 -43 391 1 gnd
rlabel metal1 68 462 68 462 7 s1
rlabel metal1 -42 314 -42 314 1 vdd
rlabel metal1 -43 218 -43 218 1 gnd
rlabel metal1 -44 136 -44 136 1 vdd
rlabel metal1 -45 40 -45 40 1 gnd
rlabel metal1 -45 -19 -45 -19 1 vdd
rlabel metal1 -46 -115 -46 -115 1 gnd
rlabel metal2 -83 324 -83 324 1 p2
rlabel metal1 -82 255 -82 255 1 c1
rlabel metal2 -85 146 -85 146 1 p3
rlabel metal1 -84 77 -84 77 1 c2
rlabel metal2 -86 -9 -86 -9 3 p4
rlabel metal1 -85 -78 -85 -78 1 c3
rlabel metal1 65 -44 65 -44 1 s4
rlabel metal1 66 111 66 111 7 s3
rlabel metal1 68 289 68 289 7 s2
<< end >>

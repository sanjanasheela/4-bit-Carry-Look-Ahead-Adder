magic
tech scmos
timestamp 1732098341
<< nwell >>
rect 133 -243 212 -185
rect 121 -677 200 -619
rect 121 -1117 200 -1059
rect 114 -1511 193 -1453
<< ntransistor >>
rect 182 -113 184 -94
rect 212 -113 214 -94
rect 138 -147 140 -128
rect 144 -309 146 -269
rect 163 -309 165 -269
rect 198 -282 200 -262
rect 170 -547 172 -528
rect 200 -547 202 -528
rect 126 -581 128 -562
rect 132 -743 134 -703
rect 151 -743 153 -703
rect 186 -716 188 -696
rect 170 -987 172 -968
rect 200 -987 202 -968
rect 126 -1021 128 -1002
rect 132 -1183 134 -1143
rect 151 -1183 153 -1143
rect 186 -1156 188 -1136
rect 163 -1381 165 -1362
rect 193 -1381 195 -1362
rect 119 -1415 121 -1396
rect 125 -1577 127 -1537
rect 144 -1577 146 -1537
rect 179 -1550 181 -1530
<< ptransistor >>
rect 138 -105 140 -65
rect 182 -71 184 -31
rect 212 -71 214 -31
rect 144 -237 146 -197
rect 163 -237 165 -197
rect 198 -237 200 -197
rect 126 -539 128 -499
rect 170 -505 172 -465
rect 200 -505 202 -465
rect 132 -671 134 -631
rect 151 -671 153 -631
rect 186 -671 188 -631
rect 126 -979 128 -939
rect 170 -945 172 -905
rect 200 -945 202 -905
rect 132 -1111 134 -1071
rect 151 -1111 153 -1071
rect 186 -1111 188 -1071
rect 119 -1373 121 -1333
rect 163 -1339 165 -1299
rect 193 -1339 195 -1299
rect 125 -1505 127 -1465
rect 144 -1505 146 -1465
rect 179 -1505 181 -1465
<< ndiffusion >>
rect 181 -113 182 -94
rect 184 -113 185 -94
rect 211 -113 212 -94
rect 214 -113 215 -94
rect 137 -147 138 -128
rect 140 -147 141 -128
rect 143 -309 144 -269
rect 146 -309 147 -269
rect 162 -309 163 -269
rect 165 -309 166 -269
rect 197 -282 198 -262
rect 200 -282 201 -262
rect 169 -547 170 -528
rect 172 -547 173 -528
rect 199 -547 200 -528
rect 202 -547 203 -528
rect 125 -581 126 -562
rect 128 -581 129 -562
rect 131 -743 132 -703
rect 134 -743 135 -703
rect 150 -743 151 -703
rect 153 -743 154 -703
rect 185 -716 186 -696
rect 188 -716 189 -696
rect 169 -987 170 -968
rect 172 -987 173 -968
rect 199 -987 200 -968
rect 202 -987 203 -968
rect 125 -1021 126 -1002
rect 128 -1021 129 -1002
rect 131 -1183 132 -1143
rect 134 -1183 135 -1143
rect 150 -1183 151 -1143
rect 153 -1183 154 -1143
rect 185 -1156 186 -1136
rect 188 -1156 189 -1136
rect 162 -1381 163 -1362
rect 165 -1381 166 -1362
rect 192 -1381 193 -1362
rect 195 -1381 196 -1362
rect 118 -1415 119 -1396
rect 121 -1415 122 -1396
rect 124 -1577 125 -1537
rect 127 -1577 128 -1537
rect 143 -1577 144 -1537
rect 146 -1577 147 -1537
rect 178 -1550 179 -1530
rect 181 -1550 182 -1530
<< pdiffusion >>
rect 137 -105 138 -65
rect 140 -105 141 -65
rect 181 -71 182 -31
rect 184 -71 185 -31
rect 211 -71 212 -31
rect 214 -71 215 -31
rect 143 -237 144 -197
rect 146 -237 147 -197
rect 162 -237 163 -197
rect 165 -237 166 -197
rect 197 -237 198 -197
rect 200 -237 201 -197
rect 125 -539 126 -499
rect 128 -539 129 -499
rect 169 -505 170 -465
rect 172 -505 173 -465
rect 199 -505 200 -465
rect 202 -505 203 -465
rect 131 -671 132 -631
rect 134 -671 135 -631
rect 150 -671 151 -631
rect 153 -671 154 -631
rect 185 -671 186 -631
rect 188 -671 189 -631
rect 125 -979 126 -939
rect 128 -979 129 -939
rect 169 -945 170 -905
rect 172 -945 173 -905
rect 199 -945 200 -905
rect 202 -945 203 -905
rect 131 -1111 132 -1071
rect 134 -1111 135 -1071
rect 150 -1111 151 -1071
rect 153 -1111 154 -1071
rect 185 -1111 186 -1071
rect 188 -1111 189 -1071
rect 118 -1373 119 -1333
rect 121 -1373 122 -1333
rect 162 -1339 163 -1299
rect 165 -1339 166 -1299
rect 192 -1339 193 -1299
rect 195 -1339 196 -1299
rect 124 -1505 125 -1465
rect 127 -1505 128 -1465
rect 143 -1505 144 -1465
rect 146 -1505 147 -1465
rect 178 -1505 179 -1465
rect 181 -1505 182 -1465
<< ndcontact >>
rect 177 -113 181 -94
rect 185 -113 189 -94
rect 207 -113 211 -94
rect 215 -113 219 -94
rect 133 -147 137 -128
rect 141 -147 145 -128
rect 139 -309 143 -269
rect 147 -309 151 -269
rect 158 -309 162 -269
rect 166 -309 170 -269
rect 193 -282 197 -262
rect 201 -282 205 -262
rect 165 -547 169 -528
rect 173 -547 177 -528
rect 195 -547 199 -528
rect 203 -547 207 -528
rect 121 -581 125 -562
rect 129 -581 133 -562
rect 127 -743 131 -703
rect 135 -743 139 -703
rect 146 -743 150 -703
rect 154 -743 158 -703
rect 181 -716 185 -696
rect 189 -716 193 -696
rect 165 -987 169 -968
rect 173 -987 177 -968
rect 195 -987 199 -968
rect 203 -987 207 -968
rect 121 -1021 125 -1002
rect 129 -1021 133 -1002
rect 127 -1183 131 -1143
rect 135 -1183 139 -1143
rect 146 -1183 150 -1143
rect 154 -1183 158 -1143
rect 181 -1156 185 -1136
rect 189 -1156 193 -1136
rect 158 -1381 162 -1362
rect 166 -1381 170 -1362
rect 188 -1381 192 -1362
rect 196 -1381 200 -1362
rect 114 -1415 118 -1396
rect 122 -1415 126 -1396
rect 120 -1577 124 -1537
rect 128 -1577 132 -1537
rect 139 -1577 143 -1537
rect 147 -1577 151 -1537
rect 174 -1550 178 -1530
rect 182 -1550 186 -1530
<< pdcontact >>
rect 133 -105 137 -65
rect 141 -105 145 -65
rect 177 -71 181 -31
rect 185 -71 189 -31
rect 207 -71 211 -31
rect 215 -71 219 -31
rect 139 -237 143 -197
rect 147 -237 151 -197
rect 158 -237 162 -197
rect 166 -237 170 -197
rect 193 -237 197 -197
rect 201 -237 205 -197
rect 121 -539 125 -499
rect 129 -539 133 -499
rect 165 -505 169 -465
rect 173 -505 177 -465
rect 195 -505 199 -465
rect 203 -505 207 -465
rect 127 -671 131 -631
rect 135 -671 139 -631
rect 146 -671 150 -631
rect 154 -671 158 -631
rect 181 -671 185 -631
rect 189 -671 193 -631
rect 121 -979 125 -939
rect 129 -979 133 -939
rect 165 -945 169 -905
rect 173 -945 177 -905
rect 195 -945 199 -905
rect 203 -945 207 -905
rect 127 -1111 131 -1071
rect 135 -1111 139 -1071
rect 146 -1111 150 -1071
rect 154 -1111 158 -1071
rect 181 -1111 185 -1071
rect 189 -1111 193 -1071
rect 114 -1373 118 -1333
rect 122 -1373 126 -1333
rect 158 -1339 162 -1299
rect 166 -1339 170 -1299
rect 188 -1339 192 -1299
rect 196 -1339 200 -1299
rect 120 -1505 124 -1465
rect 128 -1505 132 -1465
rect 139 -1505 143 -1465
rect 147 -1505 151 -1465
rect 174 -1505 178 -1465
rect 182 -1505 186 -1465
<< polysilicon >>
rect 182 -31 184 -24
rect 212 -31 214 -28
rect 138 -65 140 -62
rect 182 -74 184 -71
rect 182 -94 184 -91
rect 212 -94 214 -71
rect 138 -128 140 -105
rect 182 -120 184 -113
rect 212 -117 214 -113
rect 138 -151 140 -147
rect 144 -197 146 -194
rect 163 -197 165 -194
rect 198 -197 200 -194
rect 144 -269 146 -237
rect 163 -269 165 -237
rect 198 -262 200 -237
rect 198 -286 200 -282
rect 144 -313 146 -309
rect 163 -313 165 -309
rect 170 -465 172 -458
rect 200 -465 202 -462
rect 126 -499 128 -496
rect 170 -508 172 -505
rect 170 -528 172 -525
rect 200 -528 202 -505
rect 126 -562 128 -539
rect 170 -554 172 -547
rect 200 -551 202 -547
rect 126 -585 128 -581
rect 132 -631 134 -628
rect 151 -631 153 -628
rect 186 -631 188 -628
rect 132 -703 134 -671
rect 151 -703 153 -671
rect 186 -696 188 -671
rect 186 -720 188 -716
rect 132 -747 134 -743
rect 151 -747 153 -743
rect 170 -905 172 -898
rect 200 -905 202 -902
rect 126 -939 128 -936
rect 170 -948 172 -945
rect 170 -968 172 -965
rect 200 -968 202 -945
rect 126 -1002 128 -979
rect 170 -994 172 -987
rect 200 -991 202 -987
rect 126 -1025 128 -1021
rect 132 -1071 134 -1068
rect 151 -1071 153 -1068
rect 186 -1071 188 -1068
rect 132 -1143 134 -1111
rect 151 -1143 153 -1111
rect 186 -1136 188 -1111
rect 186 -1160 188 -1156
rect 132 -1187 134 -1183
rect 151 -1187 153 -1183
rect 163 -1299 165 -1292
rect 193 -1299 195 -1296
rect 119 -1333 121 -1330
rect 163 -1342 165 -1339
rect 163 -1362 165 -1359
rect 193 -1362 195 -1339
rect 119 -1396 121 -1373
rect 163 -1388 165 -1381
rect 193 -1385 195 -1381
rect 119 -1419 121 -1415
rect 125 -1465 127 -1462
rect 144 -1465 146 -1462
rect 179 -1465 181 -1462
rect 125 -1537 127 -1505
rect 144 -1537 146 -1505
rect 179 -1530 181 -1505
rect 179 -1554 181 -1550
rect 125 -1581 127 -1577
rect 144 -1581 146 -1577
<< polycontact >>
rect 178 -28 182 -24
rect 208 -86 212 -82
rect 134 -120 138 -116
rect 178 -120 182 -116
rect 140 -248 144 -244
rect 159 -258 163 -254
rect 194 -248 198 -244
rect 166 -462 170 -458
rect 196 -520 200 -516
rect 122 -554 126 -550
rect 166 -554 170 -550
rect 128 -682 132 -678
rect 147 -692 151 -688
rect 182 -682 186 -678
rect 166 -902 170 -898
rect 196 -960 200 -956
rect 122 -994 126 -990
rect 166 -994 170 -990
rect 128 -1122 132 -1118
rect 147 -1132 151 -1128
rect 182 -1122 186 -1118
rect 159 -1296 163 -1292
rect 189 -1354 193 -1350
rect 115 -1388 119 -1384
rect 159 -1388 163 -1384
rect 121 -1516 125 -1512
rect 140 -1526 144 -1522
rect 175 -1516 179 -1512
<< metal1 >>
rect 158 -21 211 -16
rect 158 -24 163 -21
rect 119 -28 178 -24
rect 119 -116 124 -28
rect 207 -31 211 -21
rect 130 -60 147 -56
rect 133 -65 137 -60
rect 158 -82 163 -51
rect 177 -82 181 -71
rect 185 -72 189 -71
rect 215 -81 219 -71
rect 158 -86 208 -82
rect 215 -86 224 -81
rect 229 -82 272 -81
rect 229 -86 273 -82
rect 141 -116 145 -105
rect 177 -94 181 -86
rect 215 -94 219 -86
rect 97 -120 134 -116
rect 141 -120 178 -116
rect 97 -254 100 -120
rect 141 -128 145 -120
rect 165 -123 169 -120
rect 207 -123 211 -113
rect 165 -128 211 -123
rect 133 -153 137 -147
rect 128 -157 147 -153
rect 133 -190 212 -185
rect 139 -197 143 -190
rect 158 -197 162 -190
rect 193 -197 197 -190
rect 147 -244 151 -237
rect 166 -244 170 -237
rect 201 -244 205 -237
rect 126 -248 140 -244
rect 152 -248 194 -244
rect 201 -248 267 -244
rect 201 -254 205 -248
rect 97 -258 159 -254
rect 193 -258 205 -254
rect 139 -266 147 -263
rect 193 -262 197 -258
rect 139 -269 143 -266
rect 147 -315 151 -309
rect 158 -315 162 -309
rect 147 -318 162 -315
rect 166 -321 170 -309
rect 201 -321 205 -282
rect 127 -326 211 -321
rect 146 -455 199 -450
rect 146 -458 151 -455
rect 107 -462 166 -458
rect 107 -550 112 -462
rect 195 -465 199 -455
rect 118 -494 135 -490
rect 121 -499 125 -494
rect 146 -516 151 -485
rect 165 -516 169 -505
rect 173 -506 177 -505
rect 203 -515 207 -505
rect 146 -520 196 -516
rect 203 -520 212 -515
rect 217 -516 260 -515
rect 217 -520 261 -516
rect 129 -550 133 -539
rect 165 -528 169 -520
rect 203 -528 207 -520
rect 85 -554 122 -550
rect 129 -554 166 -550
rect 85 -688 88 -554
rect 129 -562 133 -554
rect 153 -557 157 -554
rect 195 -557 199 -547
rect 153 -562 199 -557
rect 121 -587 125 -581
rect 116 -591 135 -587
rect 121 -624 200 -619
rect 127 -631 131 -624
rect 146 -631 150 -624
rect 181 -631 185 -624
rect 135 -678 139 -671
rect 154 -678 158 -671
rect 189 -678 193 -671
rect 114 -682 128 -678
rect 140 -682 182 -678
rect 189 -682 255 -678
rect 189 -688 193 -682
rect 85 -692 147 -688
rect 181 -692 193 -688
rect 127 -700 135 -697
rect 181 -696 185 -692
rect 127 -703 131 -700
rect 135 -749 139 -743
rect 146 -749 150 -743
rect 135 -752 150 -749
rect 154 -755 158 -743
rect 189 -755 193 -716
rect 115 -760 199 -755
rect 146 -895 199 -890
rect 146 -898 151 -895
rect 107 -902 166 -898
rect 107 -990 112 -902
rect 195 -905 199 -895
rect 118 -934 135 -930
rect 121 -939 125 -934
rect 146 -956 151 -925
rect 165 -956 169 -945
rect 173 -946 177 -945
rect 203 -955 207 -945
rect 146 -960 196 -956
rect 203 -960 212 -955
rect 217 -956 260 -955
rect 217 -960 261 -956
rect 129 -990 133 -979
rect 165 -968 169 -960
rect 203 -968 207 -960
rect 85 -994 122 -990
rect 129 -994 166 -990
rect 85 -1128 88 -994
rect 129 -1002 133 -994
rect 153 -997 157 -994
rect 195 -997 199 -987
rect 153 -1002 199 -997
rect 121 -1027 125 -1021
rect 116 -1031 135 -1027
rect 121 -1064 200 -1059
rect 127 -1071 131 -1064
rect 146 -1071 150 -1064
rect 181 -1071 185 -1064
rect 135 -1118 139 -1111
rect 154 -1118 158 -1111
rect 189 -1118 193 -1111
rect 114 -1122 128 -1118
rect 140 -1122 182 -1118
rect 189 -1122 255 -1118
rect 189 -1128 193 -1122
rect 85 -1132 147 -1128
rect 181 -1132 193 -1128
rect 127 -1140 135 -1137
rect 181 -1136 185 -1132
rect 127 -1143 131 -1140
rect 135 -1189 139 -1183
rect 146 -1189 150 -1183
rect 135 -1192 150 -1189
rect 154 -1195 158 -1183
rect 189 -1195 193 -1156
rect 115 -1200 199 -1195
rect 139 -1289 192 -1284
rect 139 -1292 144 -1289
rect 100 -1296 159 -1292
rect 100 -1384 105 -1296
rect 188 -1299 192 -1289
rect 111 -1328 128 -1324
rect 114 -1333 118 -1328
rect 139 -1350 144 -1319
rect 158 -1350 162 -1339
rect 166 -1340 170 -1339
rect 196 -1349 200 -1339
rect 139 -1354 189 -1350
rect 196 -1354 205 -1349
rect 210 -1350 253 -1349
rect 210 -1354 254 -1350
rect 122 -1384 126 -1373
rect 158 -1362 162 -1354
rect 196 -1362 200 -1354
rect 78 -1388 115 -1384
rect 122 -1388 159 -1384
rect 78 -1522 81 -1388
rect 122 -1396 126 -1388
rect 146 -1391 150 -1388
rect 188 -1391 192 -1381
rect 146 -1396 192 -1391
rect 114 -1421 118 -1415
rect 109 -1425 128 -1421
rect 114 -1458 193 -1453
rect 120 -1465 124 -1458
rect 139 -1465 143 -1458
rect 174 -1465 178 -1458
rect 128 -1512 132 -1505
rect 147 -1512 151 -1505
rect 182 -1512 186 -1505
rect 107 -1516 121 -1512
rect 133 -1516 175 -1512
rect 182 -1516 248 -1512
rect 182 -1522 186 -1516
rect 78 -1526 140 -1522
rect 174 -1526 186 -1522
rect 120 -1534 128 -1531
rect 174 -1530 178 -1526
rect 120 -1537 124 -1534
rect 128 -1583 132 -1577
rect 139 -1583 143 -1577
rect 128 -1586 143 -1583
rect 147 -1589 151 -1577
rect 182 -1589 186 -1550
rect 108 -1594 192 -1589
<< metal2 >>
rect 195 -13 229 -9
rect 78 -51 158 -46
rect 78 -244 82 -51
rect 195 -72 200 -13
rect 225 -17 229 -13
rect 190 -77 200 -72
rect 185 -89 190 -77
rect 224 -81 229 -17
rect 78 -249 121 -244
rect 147 -261 152 -249
rect 183 -447 217 -443
rect 66 -485 146 -480
rect 66 -678 70 -485
rect 183 -506 188 -447
rect 213 -451 217 -447
rect 178 -511 188 -506
rect 173 -523 178 -511
rect 212 -515 217 -451
rect 66 -683 109 -678
rect 135 -695 140 -683
rect 183 -887 217 -883
rect 66 -925 146 -920
rect 66 -1118 70 -925
rect 183 -946 188 -887
rect 213 -891 217 -887
rect 178 -951 188 -946
rect 173 -963 178 -951
rect 212 -955 217 -891
rect 66 -1123 109 -1118
rect 135 -1135 140 -1123
rect 176 -1281 210 -1277
rect 59 -1319 139 -1314
rect 59 -1512 63 -1319
rect 176 -1340 181 -1281
rect 206 -1285 210 -1281
rect 171 -1345 181 -1340
rect 166 -1357 171 -1345
rect 205 -1349 210 -1285
rect 59 -1517 102 -1512
rect 128 -1529 133 -1517
<< m123contact >>
rect 158 -51 163 -46
rect 185 -77 190 -72
rect 224 -86 229 -81
rect 185 -94 190 -89
rect 121 -249 126 -244
rect 147 -249 152 -244
rect 147 -266 152 -261
rect 146 -485 151 -480
rect 173 -511 178 -506
rect 212 -520 217 -515
rect 173 -528 178 -523
rect 109 -683 114 -678
rect 135 -683 140 -678
rect 135 -700 140 -695
rect 146 -925 151 -920
rect 173 -951 178 -946
rect 212 -960 217 -955
rect 173 -968 178 -963
rect 109 -1123 114 -1118
rect 135 -1123 140 -1118
rect 135 -1140 140 -1135
rect 139 -1319 144 -1314
rect 166 -1345 171 -1340
rect 205 -1354 210 -1349
rect 166 -1362 171 -1357
rect 102 -1517 107 -1512
rect 128 -1517 133 -1512
rect 128 -1534 133 -1529
<< labels >>
rlabel metal2 109 -49 109 -49 1 a1
rlabel metal1 108 -118 108 -118 1 b1
rlabel metal1 138 -58 138 -58 1 vdd
rlabel metal1 141 -156 141 -156 1 gnd
rlabel metal1 150 -189 150 -189 1 vdd
rlabel metal1 156 -324 156 -324 1 gnd
rlabel metal1 215 -247 215 -247 1 g1
rlabel metal1 237 -84 237 -84 1 p1
rlabel metal1 126 -492 126 -492 1 vdd
rlabel metal1 129 -590 129 -590 1 gnd
rlabel metal1 138 -623 138 -623 1 vdd
rlabel metal1 144 -758 144 -758 1 gnd
rlabel metal1 126 -932 126 -932 1 vdd
rlabel metal1 129 -1030 129 -1030 1 gnd
rlabel metal1 138 -1063 138 -1063 1 vdd
rlabel metal1 144 -1198 144 -1198 1 gnd
rlabel metal1 119 -1326 119 -1326 1 vdd
rlabel metal1 122 -1424 122 -1424 1 gnd
rlabel metal1 131 -1457 131 -1457 1 vdd
rlabel metal1 137 -1592 137 -1592 1 gnd
rlabel metal2 97 -483 97 -483 1 a2
rlabel metal1 96 -552 96 -552 1 b2
rlabel metal2 97 -923 97 -923 1 a3
rlabel metal1 96 -992 96 -992 1 b3
rlabel metal2 90 -1317 90 -1317 1 a4
rlabel metal1 89 -1386 89 -1386 1 b4
rlabel metal1 196 -1515 196 -1515 1 g4
rlabel metal1 218 -1352 218 -1352 1 p4
rlabel metal1 203 -1121 203 -1121 1 g3
rlabel metal1 225 -958 225 -958 1 p3
rlabel metal1 203 -681 203 -681 1 g2
rlabel metal1 225 -518 225 -518 1 p2
<< end >>
